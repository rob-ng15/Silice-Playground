`define DE10NANO 1

module SdramVga(
    input clk,
    output reg[7:0] led,

    // SDRAM
    output reg SDRAM_CLK,
    output reg SDRAM_CKE,
    output reg SDRAM_DQML,
    output reg SDRAM_DQMH,
    output reg SDRAM_nCS,
    output reg SDRAM_nWE,
    output reg SDRAM_nCAS,
    output reg SDRAM_nRAS,
    output reg [1:0] SDRAM_BA,
    output reg [12:0] SDRAM_A,
    // inout [15:0] SDRAM_DQ,
    inout [7:0] SDRAM_DQ,

    // VGA
    output reg vga_hs,
    output reg vga_vs,
    output reg [5:0] vga_r,
    output reg [5:0] vga_g,
    output reg [5:0] vga_b,

    // uart via GPIO pins
    output tx,
    input rx,
    
    // user button and switches
    input   BUTTON0,
    input   BUTTON1,
    input   SWITCH0,
    input   SWITCH1,
    input   SWITCH2,
    input   SWITCH3    
);

wire [7:0]  __main_out_led;

wire        __main_out_sdram_clk;
wire        __main_out_sdram_cle;
wire        __main_out_sdram_dqm;
wire        __main_out_sdram_cs;
wire        __main_out_sdram_we;
wire        __main_out_sdram_cas;
wire        __main_out_sdram_ras;
wire [1:0]  __main_out_sdram_ba;
wire [12:0] __main_out_sdram_a;
  
wire        __main_out_vga_hs;
wire        __main_out_vga_vs;
wire [5:0]  __main_out_vga_r;
wire [5:0]  __main_out_vga_g;
wire [5:0]  __main_out_vga_b;

reg [31:0] RST_d;
reg [31:0] RST_q;

reg ready = 0;

always @* begin
  RST_d = RST_q >> 1;
end

always @(posedge clk) begin
  if (ready) begin
    RST_q <= RST_d;
  end else begin
    ready <= 1;
    RST_q <= 32'b111111111111111111111111111111;
  end
end

wire reset_main;
assign reset_main = RST_q[0];
wire run_main;
assign run_main = 1'b1;

// Create 1hz (1 second counter)
reg [31:0] counter50mhz;
reg [15:0] counter1hz;
always @(posedge clk) begin
    if( counter50mhz == 50000000 ) begin
        counter1hz <= counter1hz + 1;
        counter50mhz <= 0;
    end else begin
        counter50mhz <= counter50mhz + 1;
    end
end 

// UART tx and rx
wire [7:0] uart_tx_data;
wire uart_tx_valid;
wire uart_tx_busy;
wire uart_tx_done;
wire [7:0] uart_rx_data;
wire uart_rx_valid;
wire uart_rx_ready;
wire uart_serial_tx;

// UART from https://github.com/cyrozap/osdvu
uart uart0(
    .clk(clk), // The master clock for this module
    .rst(reset_main), // Synchronous reset
    .rx(rx), // Incoming serial line
    .tx(tx), // Outgoing serial line
    .transmit(uart_tx_valid), // Signal to transmit
    .tx_byte(uart_tx_data), // Byte to transmit
    .received(uart_rx_valid), // Indicated that a byte has been received
    .rx_byte(uart_rx_data), // Byte received
    .is_receiving(), // Low when receive line is idle
    .is_transmitting(uart_tx_busy),// Low when transmit line is idle
    .recv_error() // Indicates error in receiving packet.
);

M_main __main(
  // CLK and RESET
  .clock(clk),
  .reset(reset_main),
  .in_run(run_main),
  
  // LEDS
  .out_led(__main_out_led),

  // BUTTONS and SWITCHES (combined)
  .in_buttons( {2'b0, SWITCH3, SWITCH2, SWITCH1, SWITCH0, BUTTON1, BUTTON0} ),
  
  .inout_sdram_dq(SDRAM_DQ[7:0]),
  .out_sdram_clk(__main_out_sdram_clk),
  .out_sdram_cle(__main_out_sdram_cle),
  .out_sdram_dqm(__main_out_sdram_dqm),
  .out_sdram_cs(__main_out_sdram_cs),
  .out_sdram_we(__main_out_sdram_we),
  .out_sdram_cas(__main_out_sdram_cas),
  .out_sdram_ras(__main_out_sdram_ras),
  .out_sdram_ba(__main_out_sdram_ba),
  .out_sdram_a(__main_out_sdram_a),
  .out_video_hs(__main_out_vga_hs),
  .out_video_vs(__main_out_vga_vs),
  .out_video_r(__main_out_vga_r),
  .out_video_g(__main_out_vga_g),
  .out_video_b(__main_out_vga_b),

  // UART
  .out_uart_tx_data( uart_tx_data ),
  .out_uart_tx_valid( uart_tx_valid ),
  .in_uart_tx_busy( uart_tx_busy ),
  .in_uart_tx_done( uart_tx_done ),

  .in_uart_rx_data( uart_rx_data ),
  .in_uart_rx_valid( uart_rx_valid ),
    
  .in_timer1hz ( counter1hz )
);

always @* begin

  led          = __main_out_led;

  SDRAM_CLK    = __main_out_sdram_clk;
  SDRAM_CKE    = __main_out_sdram_cle;
  SDRAM_DQML   = __main_out_sdram_dqm;
  SDRAM_DQMH   = 0;
  SDRAM_nCS    = __main_out_sdram_cs;
  SDRAM_nWE    = __main_out_sdram_we;
  SDRAM_nCAS   = __main_out_sdram_cas;
  SDRAM_nRAS   = __main_out_sdram_ras;
  SDRAM_BA     = __main_out_sdram_ba;
  SDRAM_A      = __main_out_sdram_a;
  vga_hs       = __main_out_vga_hs;
  vga_vs       = __main_out_vga_vs;
  vga_r        = __main_out_vga_r;
  vga_g        = __main_out_vga_g;
  vga_b        = __main_out_vga_b;

end

endmodule

`timescale 1ns/10ps

module  de10nano_clk_100_25(
	// interface 'refclk'
	input refclk,
	// interface 'reset'
	input rst,
	// interface 'outclk0'
	output outclk_0,
	// interface 'outclk1'
	output outclk_1,
	// interface 'locked'
	output locked
);

	altera_pll #(
		.fractional_vco_multiplier("true"),
		.reference_clock_frequency("50.0 MHz"),
		.operation_mode("direct"),
		.number_of_clocks(2),
		.output_clock_frequency0("100.000000 MHz"),
		.phase_shift0("0 ps"),
		.duty_cycle0(50),
		.output_clock_frequency1("25.000000 MHz"),
		.phase_shift1("0 ps"),
		.duty_cycle1(50),
		.output_clock_frequency2("0 MHz"),
		.phase_shift2("0 ps"),
		.duty_cycle2(50),
		.output_clock_frequency3("0 MHz"),
		.phase_shift3("0 ps"),
		.duty_cycle3(50),
		.output_clock_frequency4("0 MHz"),
		.phase_shift4("0 ps"),
		.duty_cycle4(50),
		.output_clock_frequency5("0 MHz"),
		.phase_shift5("0 ps"),
		.duty_cycle5(50),
		.output_clock_frequency6("0 MHz"),
		.phase_shift6("0 ps"),
		.duty_cycle6(50),
		.output_clock_frequency7("0 MHz"),
		.phase_shift7("0 ps"),
		.duty_cycle7(50),
		.output_clock_frequency8("0 MHz"),
		.phase_shift8("0 ps"),
		.duty_cycle8(50),
		.output_clock_frequency9("0 MHz"),
		.phase_shift9("0 ps"),
		.duty_cycle9(50),
		.output_clock_frequency10("0 MHz"),
		.phase_shift10("0 ps"),
		.duty_cycle10(50),
		.output_clock_frequency11("0 MHz"),
		.phase_shift11("0 ps"),
		.duty_cycle11(50),
		.output_clock_frequency12("0 MHz"),
		.phase_shift12("0 ps"),
		.duty_cycle12(50),
		.output_clock_frequency13("0 MHz"),
		.phase_shift13("0 ps"),
		.duty_cycle13(50),
		.output_clock_frequency14("0 MHz"),
		.phase_shift14("0 ps"),
		.duty_cycle14(50),
		.output_clock_frequency15("0 MHz"),
		.phase_shift15("0 ps"),
		.duty_cycle15(50),
		.output_clock_frequency16("0 MHz"),
		.phase_shift16("0 ps"),
		.duty_cycle16(50),
		.output_clock_frequency17("0 MHz"),
		.phase_shift17("0 ps"),
		.duty_cycle17(50),
		.pll_type("General"),
		.pll_subtype("General")
	) altera_pll_i (
		.rst	(rst),
		.outclk	({outclk_1, outclk_0}),
		.locked	(locked),
		.fboutclk	( ),
		.fbclk	(1'b0),
		.refclk	(refclk)
	);
endmodule



module reset_conditioner (
    input rcclk,
    input in,
    output reg out
  );  
  reg [7:0] counter_d,counter_q;
  always @* begin
    counter_d = counter_q;
    if (counter_q == 0) begin
      out = 0;
    end else begin
      out = 1;
      counter_d = counter_q + 1;
    end
  end  
  always @(posedge rcclk) begin
    if (in == 1'b1) begin
      counter_q <= 1;
    end else begin
      counter_q <= counter_d;
    end
  end 
endmodule


module M_vga (
out_vga_hs,
out_vga_vs,
out_active,
out_vblank,
out_vga_x,
out_vga_y,
in_run,
out_done,
reset,
clock
);
output  [0:0] out_vga_hs;
output  [0:0] out_vga_vs;
output  [0:0] out_active;
output  [0:0] out_vblank;
output  [9:0] out_vga_x;
output  [9:0] out_vga_y;
input in_run;
output out_done;
input reset;
input clock;
wire  [9:0] _c_H_FRT_PORCH;
assign _c_H_FRT_PORCH = 16;
wire  [9:0] _c_H_SYNCH;
assign _c_H_SYNCH = 96;
wire  [9:0] _c_H_BCK_PORCH;
assign _c_H_BCK_PORCH = 48;
wire  [9:0] _c_H_RES;
assign _c_H_RES = 640;
wire  [9:0] _c_V_FRT_PORCH;
assign _c_V_FRT_PORCH = 10;
wire  [9:0] _c_V_SYNCH;
assign _c_V_SYNCH = 2;
wire  [9:0] _c_V_BCK_PORCH;
assign _c_V_BCK_PORCH = 33;
wire  [9:0] _c_V_RES;
assign _c_V_RES = 480;
reg  [9:0] _t_HS_START;
reg  [9:0] _t_HS_END;
reg  [9:0] _t_HA_START;
reg  [9:0] _t_H_END;
reg  [9:0] _t_VS_START;
reg  [9:0] _t_VS_END;
reg  [9:0] _t_VA_START;
reg  [9:0] _t_V_END;

reg  [9:0] _d_xcount;
reg  [9:0] _q_xcount;
reg  [9:0] _d_ycount;
reg  [9:0] _q_ycount;
reg  [0:0] _d_vga_hs,_q_vga_hs;
reg  [0:0] _d_vga_vs,_q_vga_vs;
reg  [0:0] _d_active,_q_active;
reg  [0:0] _d_vblank,_q_vblank;
reg  [9:0] _d_vga_x,_q_vga_x;
reg  [9:0] _d_vga_y,_q_vga_y;
reg  [1:0] _d_index,_q_index;
assign out_vga_hs = _d_vga_hs;
assign out_vga_vs = _d_vga_vs;
assign out_active = _d_active;
assign out_vblank = _d_vblank;
assign out_vga_x = _d_vga_x;
assign out_vga_y = _d_vga_y;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_xcount <= 0;
_q_ycount <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_xcount <= _d_xcount;
_q_ycount <= _d_ycount;
_q_index <= _d_index;
  end
_q_vga_hs <= _d_vga_hs;
_q_vga_vs <= _d_vga_vs;
_q_active <= _d_active;
_q_vblank <= _d_vblank;
_q_vga_x <= _d_vga_x;
_q_vga_y <= _d_vga_y;
end




always @* begin
_d_xcount = _q_xcount;
_d_ycount = _q_ycount;
_d_vga_hs = _q_vga_hs;
_d_vga_vs = _q_vga_vs;
_d_active = _q_active;
_d_vblank = _q_vblank;
_d_vga_x = _q_vga_x;
_d_vga_y = _q_vga_y;
_d_index = _q_index;
_t_HS_START = 0;
_t_HS_END = 0;
_t_HA_START = 0;
_t_H_END = 0;
_t_VS_START = 0;
_t_VS_END = 0;
_t_VA_START = 0;
_t_V_END = 0;
// _always_pre
_t_HS_START = _c_H_FRT_PORCH;
_t_HS_END = _c_H_FRT_PORCH+_c_H_SYNCH;
_t_HA_START = _c_H_FRT_PORCH+_c_H_SYNCH+_c_H_BCK_PORCH;
_t_H_END = _c_H_FRT_PORCH+_c_H_SYNCH+_c_H_BCK_PORCH+_c_H_RES;
_t_VS_START = _c_V_FRT_PORCH;
_t_VS_END = _c_V_FRT_PORCH+_c_V_SYNCH;
_t_VA_START = _c_V_FRT_PORCH+_c_V_SYNCH+_c_V_BCK_PORCH;
_t_V_END = _c_V_FRT_PORCH+_c_V_SYNCH+_c_V_BCK_PORCH+_c_V_RES;
_d_vga_hs = ~((_q_xcount>=_t_HS_START&&_q_xcount<_t_HS_END));
_d_vga_vs = ~((_q_ycount>=_t_VS_START&&_q_ycount<_t_VS_END));
_d_active = (_q_xcount>=_t_HA_START&&_q_xcount<_t_H_END)&&(_q_ycount>=_t_VA_START&&_q_ycount<_t_V_END);
_d_vblank = (_q_ycount<_t_VA_START);
_d_index = 3;
case (_q_index)
0: begin
// _top
// var inits
_t_HS_START = 0;
_t_HS_END = 0;
_t_HA_START = 0;
_t_H_END = 0;
_t_VS_START = 0;
_t_VS_END = 0;
_t_VA_START = 0;
_t_V_END = 0;
_d_xcount = 0;
_d_ycount = 0;
// --
_d_xcount = 0;
_d_ycount = 0;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (_d_active) begin
// __block_5
// __block_7
_d_vga_x = _q_xcount-_t_HA_START;
_d_vga_y = _q_ycount-_t_VA_START;
// __block_8
end else begin
// __block_6
end
// __block_9
if (_q_xcount==_t_H_END-1) begin
// __block_10
// __block_12
_d_xcount = 0;
if (_q_ycount==_t_V_END-1) begin
// __block_13
// __block_15
_d_ycount = 0;
// __block_16
end else begin
// __block_14
// __block_17
_d_ycount = _q_ycount+1;
// __block_18
end
// __block_19
// __block_20
end else begin
// __block_11
// __block_21
_d_xcount = _q_xcount+1;
// __block_22
end
// __block_23
// __block_24
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of vga
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_multiplex_display_mem_character(
input      [0:0]             in_character_wenable0,
input       [7:0]     in_character_wdata0,
input      [11:0]                in_character_addr0,
input      [0:0]             in_character_wenable1,
input      [7:0]                 in_character_wdata1,
input      [11:0]                in_character_addr1,
output reg  [7:0]     out_character_rdata0,
output reg  [7:0]     out_character_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2399:0];
always @(posedge clock0) begin
  if (in_character_wenable0) begin
    buffer[in_character_addr0] <= in_character_wdata0;
  end else begin
    out_character_rdata0 <= buffer[in_character_addr0];
  end
end
always @(posedge clock1) begin
  if (in_character_wenable1) begin
    buffer[in_character_addr1] <= in_character_wdata1;
  end else begin
    out_character_rdata1 <= buffer[in_character_addr1];
  end
end
initial begin
 buffer[0] = 0;
 buffer[1] = 1;
 buffer[2] = 2;
 buffer[3] = 3;
 buffer[4] = 4;
 buffer[5] = 5;
 buffer[6] = 6;
 buffer[7] = 7;
 buffer[8] = 8;
 buffer[9] = 9;
 buffer[10] = 10;
 buffer[11] = 11;
 buffer[12] = 12;
 buffer[13] = 13;
 buffer[14] = 14;
 buffer[15] = 15;
 buffer[16] = 16;
 buffer[17] = 17;
 buffer[18] = 18;
 buffer[19] = 19;
 buffer[20] = 20;
 buffer[21] = 21;
 buffer[22] = 22;
 buffer[23] = 23;
 buffer[24] = 24;
 buffer[25] = 25;
 buffer[26] = 26;
 buffer[27] = 27;
 buffer[28] = 28;
 buffer[29] = 29;
 buffer[30] = 30;
 buffer[31] = 31;
 buffer[32] = 32;
 buffer[33] = 33;
 buffer[34] = 34;
 buffer[35] = 35;
 buffer[36] = 36;
 buffer[37] = 37;
 buffer[38] = 38;
 buffer[39] = 39;
 buffer[40] = 40;
 buffer[41] = 41;
 buffer[42] = 42;
 buffer[43] = 43;
 buffer[44] = 44;
 buffer[45] = 45;
 buffer[46] = 46;
 buffer[47] = 47;
 buffer[48] = 48;
 buffer[49] = 49;
 buffer[50] = 50;
 buffer[51] = 51;
 buffer[52] = 52;
 buffer[53] = 53;
 buffer[54] = 54;
 buffer[55] = 55;
 buffer[56] = 56;
 buffer[57] = 57;
 buffer[58] = 58;
 buffer[59] = 59;
 buffer[60] = 60;
 buffer[61] = 61;
 buffer[62] = 62;
 buffer[63] = 63;
 buffer[64] = 64;
 buffer[65] = 65;
 buffer[66] = 66;
 buffer[67] = 67;
 buffer[68] = 68;
 buffer[69] = 69;
 buffer[70] = 70;
 buffer[71] = 71;
 buffer[72] = 72;
 buffer[73] = 73;
 buffer[74] = 74;
 buffer[75] = 75;
 buffer[76] = 76;
 buffer[77] = 77;
 buffer[78] = 78;
 buffer[79] = 79;
 buffer[80] = 80;
 buffer[81] = 81;
 buffer[82] = 82;
 buffer[83] = 83;
 buffer[84] = 84;
 buffer[85] = 85;
 buffer[86] = 86;
 buffer[87] = 87;
 buffer[88] = 88;
 buffer[89] = 89;
 buffer[90] = 90;
 buffer[91] = 91;
 buffer[92] = 92;
 buffer[93] = 93;
 buffer[94] = 94;
 buffer[95] = 95;
 buffer[96] = 96;
 buffer[97] = 97;
 buffer[98] = 98;
 buffer[99] = 99;
 buffer[100] = 100;
 buffer[101] = 101;
 buffer[102] = 102;
 buffer[103] = 103;
 buffer[104] = 104;
 buffer[105] = 105;
 buffer[106] = 106;
 buffer[107] = 107;
 buffer[108] = 108;
 buffer[109] = 109;
 buffer[110] = 110;
 buffer[111] = 111;
 buffer[112] = 112;
 buffer[113] = 113;
 buffer[114] = 114;
 buffer[115] = 115;
 buffer[116] = 116;
 buffer[117] = 117;
 buffer[118] = 118;
 buffer[119] = 119;
 buffer[120] = 120;
 buffer[121] = 121;
 buffer[122] = 122;
 buffer[123] = 123;
 buffer[124] = 124;
 buffer[125] = 125;
 buffer[126] = 126;
 buffer[127] = 127;
 buffer[128] = 128;
 buffer[129] = 129;
 buffer[130] = 130;
 buffer[131] = 131;
 buffer[132] = 132;
 buffer[133] = 133;
 buffer[134] = 134;
 buffer[135] = 135;
 buffer[136] = 136;
 buffer[137] = 137;
 buffer[138] = 138;
 buffer[139] = 139;
 buffer[140] = 140;
 buffer[141] = 141;
 buffer[142] = 142;
 buffer[143] = 143;
 buffer[144] = 144;
 buffer[145] = 145;
 buffer[146] = 146;
 buffer[147] = 147;
 buffer[148] = 148;
 buffer[149] = 149;
 buffer[150] = 150;
 buffer[151] = 151;
 buffer[152] = 152;
 buffer[153] = 153;
 buffer[154] = 154;
 buffer[155] = 155;
 buffer[156] = 156;
 buffer[157] = 157;
 buffer[158] = 158;
 buffer[159] = 159;
 buffer[160] = 160;
 buffer[161] = 161;
 buffer[162] = 162;
 buffer[163] = 163;
 buffer[164] = 164;
 buffer[165] = 165;
 buffer[166] = 166;
 buffer[167] = 167;
 buffer[168] = 168;
 buffer[169] = 169;
 buffer[170] = 170;
 buffer[171] = 171;
 buffer[172] = 172;
 buffer[173] = 173;
 buffer[174] = 174;
 buffer[175] = 175;
 buffer[176] = 176;
 buffer[177] = 177;
 buffer[178] = 178;
 buffer[179] = 179;
 buffer[180] = 180;
 buffer[181] = 181;
 buffer[182] = 182;
 buffer[183] = 183;
 buffer[184] = 184;
 buffer[185] = 185;
 buffer[186] = 186;
 buffer[187] = 187;
 buffer[188] = 188;
 buffer[189] = 189;
 buffer[190] = 190;
 buffer[191] = 191;
 buffer[192] = 192;
 buffer[193] = 193;
 buffer[194] = 194;
 buffer[195] = 195;
 buffer[196] = 196;
 buffer[197] = 197;
 buffer[198] = 198;
 buffer[199] = 199;
 buffer[200] = 200;
 buffer[201] = 201;
 buffer[202] = 202;
 buffer[203] = 203;
 buffer[204] = 204;
 buffer[205] = 205;
 buffer[206] = 206;
 buffer[207] = 207;
 buffer[208] = 208;
 buffer[209] = 209;
 buffer[210] = 210;
 buffer[211] = 211;
 buffer[212] = 212;
 buffer[213] = 213;
 buffer[214] = 214;
 buffer[215] = 215;
 buffer[216] = 216;
 buffer[217] = 217;
 buffer[218] = 218;
 buffer[219] = 219;
 buffer[220] = 220;
 buffer[221] = 221;
 buffer[222] = 222;
 buffer[223] = 223;
 buffer[224] = 224;
 buffer[225] = 225;
 buffer[226] = 226;
 buffer[227] = 227;
 buffer[228] = 228;
 buffer[229] = 229;
 buffer[230] = 230;
 buffer[231] = 231;
 buffer[232] = 232;
 buffer[233] = 233;
 buffer[234] = 234;
 buffer[235] = 235;
 buffer[236] = 236;
 buffer[237] = 237;
 buffer[238] = 238;
 buffer[239] = 239;
 buffer[240] = 240;
 buffer[241] = 241;
 buffer[242] = 242;
 buffer[243] = 243;
 buffer[244] = 244;
 buffer[245] = 245;
 buffer[246] = 246;
 buffer[247] = 247;
 buffer[248] = 248;
 buffer[249] = 249;
 buffer[250] = 250;
 buffer[251] = 251;
 buffer[252] = 252;
 buffer[253] = 253;
 buffer[254] = 254;
 buffer[255] = 255;
 buffer[256] = 256;
 buffer[257] = 257;
 buffer[258] = 258;
 buffer[259] = 259;
 buffer[260] = 260;
 buffer[261] = 261;
 buffer[262] = 262;
 buffer[263] = 263;
 buffer[264] = 264;
 buffer[265] = 265;
 buffer[266] = 266;
 buffer[267] = 267;
 buffer[268] = 268;
 buffer[269] = 269;
 buffer[270] = 270;
 buffer[271] = 271;
 buffer[272] = 272;
 buffer[273] = 273;
 buffer[274] = 274;
 buffer[275] = 275;
 buffer[276] = 276;
 buffer[277] = 277;
 buffer[278] = 278;
 buffer[279] = 279;
 buffer[280] = 280;
 buffer[281] = 281;
 buffer[282] = 282;
 buffer[283] = 283;
 buffer[284] = 284;
 buffer[285] = 285;
 buffer[286] = 286;
 buffer[287] = 287;
 buffer[288] = 288;
 buffer[289] = 289;
 buffer[290] = 290;
 buffer[291] = 291;
 buffer[292] = 292;
 buffer[293] = 293;
 buffer[294] = 294;
 buffer[295] = 295;
 buffer[296] = 296;
 buffer[297] = 297;
 buffer[298] = 298;
 buffer[299] = 299;
 buffer[300] = 300;
 buffer[301] = 301;
 buffer[302] = 302;
 buffer[303] = 303;
 buffer[304] = 304;
 buffer[305] = 305;
 buffer[306] = 306;
 buffer[307] = 307;
 buffer[308] = 308;
 buffer[309] = 309;
 buffer[310] = 310;
 buffer[311] = 311;
 buffer[312] = 312;
 buffer[313] = 313;
 buffer[314] = 314;
 buffer[315] = 315;
 buffer[316] = 316;
 buffer[317] = 317;
 buffer[318] = 318;
 buffer[319] = 319;
 buffer[320] = 320;
 buffer[321] = 321;
 buffer[322] = 322;
 buffer[323] = 323;
 buffer[324] = 324;
 buffer[325] = 325;
 buffer[326] = 326;
 buffer[327] = 327;
 buffer[328] = 328;
 buffer[329] = 329;
 buffer[330] = 330;
 buffer[331] = 331;
 buffer[332] = 332;
 buffer[333] = 333;
 buffer[334] = 334;
 buffer[335] = 335;
 buffer[336] = 336;
 buffer[337] = 337;
 buffer[338] = 338;
 buffer[339] = 339;
 buffer[340] = 340;
 buffer[341] = 341;
 buffer[342] = 342;
 buffer[343] = 343;
 buffer[344] = 344;
 buffer[345] = 345;
 buffer[346] = 346;
 buffer[347] = 347;
 buffer[348] = 348;
 buffer[349] = 349;
 buffer[350] = 350;
 buffer[351] = 351;
 buffer[352] = 352;
 buffer[353] = 353;
 buffer[354] = 354;
 buffer[355] = 355;
 buffer[356] = 356;
 buffer[357] = 357;
 buffer[358] = 358;
 buffer[359] = 359;
 buffer[360] = 360;
 buffer[361] = 361;
 buffer[362] = 362;
 buffer[363] = 363;
 buffer[364] = 364;
 buffer[365] = 365;
 buffer[366] = 366;
 buffer[367] = 367;
 buffer[368] = 368;
 buffer[369] = 369;
 buffer[370] = 370;
 buffer[371] = 371;
 buffer[372] = 372;
 buffer[373] = 373;
 buffer[374] = 374;
 buffer[375] = 375;
 buffer[376] = 376;
 buffer[377] = 377;
 buffer[378] = 378;
 buffer[379] = 379;
 buffer[380] = 380;
 buffer[381] = 381;
 buffer[382] = 382;
 buffer[383] = 383;
 buffer[384] = 384;
 buffer[385] = 385;
 buffer[386] = 386;
 buffer[387] = 387;
 buffer[388] = 388;
 buffer[389] = 389;
 buffer[390] = 390;
 buffer[391] = 391;
 buffer[392] = 392;
 buffer[393] = 393;
 buffer[394] = 394;
 buffer[395] = 395;
 buffer[396] = 396;
 buffer[397] = 397;
 buffer[398] = 398;
 buffer[399] = 399;
 buffer[400] = 400;
 buffer[401] = 401;
 buffer[402] = 402;
 buffer[403] = 403;
 buffer[404] = 404;
 buffer[405] = 405;
 buffer[406] = 406;
 buffer[407] = 407;
 buffer[408] = 408;
 buffer[409] = 409;
 buffer[410] = 410;
 buffer[411] = 411;
 buffer[412] = 412;
 buffer[413] = 413;
 buffer[414] = 414;
 buffer[415] = 415;
 buffer[416] = 416;
 buffer[417] = 417;
 buffer[418] = 418;
 buffer[419] = 419;
 buffer[420] = 420;
 buffer[421] = 421;
 buffer[422] = 422;
 buffer[423] = 423;
 buffer[424] = 424;
 buffer[425] = 425;
 buffer[426] = 426;
 buffer[427] = 427;
 buffer[428] = 428;
 buffer[429] = 429;
 buffer[430] = 430;
 buffer[431] = 431;
 buffer[432] = 432;
 buffer[433] = 433;
 buffer[434] = 434;
 buffer[435] = 435;
 buffer[436] = 436;
 buffer[437] = 437;
 buffer[438] = 438;
 buffer[439] = 439;
 buffer[440] = 440;
 buffer[441] = 441;
 buffer[442] = 442;
 buffer[443] = 443;
 buffer[444] = 444;
 buffer[445] = 445;
 buffer[446] = 446;
 buffer[447] = 447;
 buffer[448] = 448;
 buffer[449] = 449;
 buffer[450] = 450;
 buffer[451] = 451;
 buffer[452] = 452;
 buffer[453] = 453;
 buffer[454] = 454;
 buffer[455] = 455;
 buffer[456] = 456;
 buffer[457] = 457;
 buffer[458] = 458;
 buffer[459] = 459;
 buffer[460] = 460;
 buffer[461] = 461;
 buffer[462] = 462;
 buffer[463] = 463;
 buffer[464] = 464;
 buffer[465] = 465;
 buffer[466] = 466;
 buffer[467] = 467;
 buffer[468] = 468;
 buffer[469] = 469;
 buffer[470] = 470;
 buffer[471] = 471;
 buffer[472] = 472;
 buffer[473] = 473;
 buffer[474] = 474;
 buffer[475] = 475;
 buffer[476] = 476;
 buffer[477] = 477;
 buffer[478] = 478;
 buffer[479] = 479;
 buffer[480] = 480;
 buffer[481] = 481;
 buffer[482] = 482;
 buffer[483] = 483;
 buffer[484] = 484;
 buffer[485] = 485;
 buffer[486] = 486;
 buffer[487] = 487;
 buffer[488] = 488;
 buffer[489] = 489;
 buffer[490] = 490;
 buffer[491] = 491;
 buffer[492] = 492;
 buffer[493] = 493;
 buffer[494] = 494;
 buffer[495] = 495;
 buffer[496] = 496;
 buffer[497] = 497;
 buffer[498] = 498;
 buffer[499] = 499;
 buffer[500] = 500;
 buffer[501] = 501;
 buffer[502] = 502;
 buffer[503] = 503;
 buffer[504] = 504;
 buffer[505] = 505;
 buffer[506] = 506;
 buffer[507] = 507;
 buffer[508] = 508;
 buffer[509] = 509;
 buffer[510] = 510;
 buffer[511] = 511;
 buffer[512] = 512;
 buffer[513] = 513;
 buffer[514] = 514;
 buffer[515] = 515;
 buffer[516] = 516;
 buffer[517] = 517;
 buffer[518] = 518;
 buffer[519] = 519;
 buffer[520] = 520;
 buffer[521] = 521;
 buffer[522] = 522;
 buffer[523] = 523;
 buffer[524] = 524;
 buffer[525] = 525;
 buffer[526] = 526;
 buffer[527] = 527;
 buffer[528] = 528;
 buffer[529] = 529;
 buffer[530] = 530;
 buffer[531] = 531;
 buffer[532] = 532;
 buffer[533] = 533;
 buffer[534] = 534;
 buffer[535] = 535;
 buffer[536] = 536;
 buffer[537] = 537;
 buffer[538] = 538;
 buffer[539] = 539;
 buffer[540] = 540;
 buffer[541] = 541;
 buffer[542] = 542;
 buffer[543] = 543;
 buffer[544] = 544;
 buffer[545] = 545;
 buffer[546] = 546;
 buffer[547] = 547;
 buffer[548] = 548;
 buffer[549] = 549;
 buffer[550] = 550;
 buffer[551] = 551;
 buffer[552] = 552;
 buffer[553] = 553;
 buffer[554] = 554;
 buffer[555] = 555;
 buffer[556] = 556;
 buffer[557] = 557;
 buffer[558] = 558;
 buffer[559] = 559;
 buffer[560] = 560;
 buffer[561] = 561;
 buffer[562] = 562;
 buffer[563] = 563;
 buffer[564] = 564;
 buffer[565] = 565;
 buffer[566] = 566;
 buffer[567] = 567;
 buffer[568] = 568;
 buffer[569] = 569;
 buffer[570] = 570;
 buffer[571] = 571;
 buffer[572] = 572;
 buffer[573] = 573;
 buffer[574] = 574;
 buffer[575] = 575;
 buffer[576] = 576;
 buffer[577] = 577;
 buffer[578] = 578;
 buffer[579] = 579;
 buffer[580] = 580;
 buffer[581] = 581;
 buffer[582] = 582;
 buffer[583] = 583;
 buffer[584] = 584;
 buffer[585] = 585;
 buffer[586] = 586;
 buffer[587] = 587;
 buffer[588] = 588;
 buffer[589] = 589;
 buffer[590] = 590;
 buffer[591] = 591;
 buffer[592] = 592;
 buffer[593] = 593;
 buffer[594] = 594;
 buffer[595] = 595;
 buffer[596] = 596;
 buffer[597] = 597;
 buffer[598] = 598;
 buffer[599] = 599;
 buffer[600] = 600;
 buffer[601] = 601;
 buffer[602] = 602;
 buffer[603] = 603;
 buffer[604] = 604;
 buffer[605] = 605;
 buffer[606] = 606;
 buffer[607] = 607;
 buffer[608] = 608;
 buffer[609] = 609;
 buffer[610] = 610;
 buffer[611] = 611;
 buffer[612] = 612;
 buffer[613] = 613;
 buffer[614] = 614;
 buffer[615] = 615;
 buffer[616] = 616;
 buffer[617] = 617;
 buffer[618] = 618;
 buffer[619] = 619;
 buffer[620] = 620;
 buffer[621] = 621;
 buffer[622] = 622;
 buffer[623] = 623;
 buffer[624] = 624;
 buffer[625] = 625;
 buffer[626] = 626;
 buffer[627] = 627;
 buffer[628] = 628;
 buffer[629] = 629;
 buffer[630] = 630;
 buffer[631] = 631;
 buffer[632] = 632;
 buffer[633] = 633;
 buffer[634] = 634;
 buffer[635] = 635;
 buffer[636] = 636;
 buffer[637] = 637;
 buffer[638] = 638;
 buffer[639] = 639;
 buffer[640] = 640;
 buffer[641] = 641;
 buffer[642] = 642;
 buffer[643] = 643;
 buffer[644] = 644;
 buffer[645] = 645;
 buffer[646] = 646;
 buffer[647] = 647;
 buffer[648] = 648;
 buffer[649] = 649;
 buffer[650] = 650;
 buffer[651] = 651;
 buffer[652] = 652;
 buffer[653] = 653;
 buffer[654] = 654;
 buffer[655] = 655;
 buffer[656] = 656;
 buffer[657] = 657;
 buffer[658] = 658;
 buffer[659] = 659;
 buffer[660] = 660;
 buffer[661] = 661;
 buffer[662] = 662;
 buffer[663] = 663;
 buffer[664] = 664;
 buffer[665] = 665;
 buffer[666] = 666;
 buffer[667] = 667;
 buffer[668] = 668;
 buffer[669] = 669;
 buffer[670] = 670;
 buffer[671] = 671;
 buffer[672] = 672;
 buffer[673] = 673;
 buffer[674] = 674;
 buffer[675] = 675;
 buffer[676] = 676;
 buffer[677] = 677;
 buffer[678] = 678;
 buffer[679] = 679;
 buffer[680] = 680;
 buffer[681] = 681;
 buffer[682] = 682;
 buffer[683] = 683;
 buffer[684] = 684;
 buffer[685] = 685;
 buffer[686] = 686;
 buffer[687] = 687;
 buffer[688] = 688;
 buffer[689] = 689;
 buffer[690] = 690;
 buffer[691] = 691;
 buffer[692] = 692;
 buffer[693] = 693;
 buffer[694] = 694;
 buffer[695] = 695;
 buffer[696] = 696;
 buffer[697] = 697;
 buffer[698] = 698;
 buffer[699] = 699;
 buffer[700] = 700;
 buffer[701] = 701;
 buffer[702] = 702;
 buffer[703] = 703;
 buffer[704] = 704;
 buffer[705] = 705;
 buffer[706] = 706;
 buffer[707] = 707;
 buffer[708] = 708;
 buffer[709] = 709;
 buffer[710] = 710;
 buffer[711] = 711;
 buffer[712] = 712;
 buffer[713] = 713;
 buffer[714] = 714;
 buffer[715] = 715;
 buffer[716] = 716;
 buffer[717] = 717;
 buffer[718] = 718;
 buffer[719] = 719;
 buffer[720] = 720;
 buffer[721] = 721;
 buffer[722] = 722;
 buffer[723] = 723;
 buffer[724] = 724;
 buffer[725] = 725;
 buffer[726] = 726;
 buffer[727] = 727;
 buffer[728] = 728;
 buffer[729] = 729;
 buffer[730] = 730;
 buffer[731] = 731;
 buffer[732] = 732;
 buffer[733] = 733;
 buffer[734] = 734;
 buffer[735] = 735;
 buffer[736] = 736;
 buffer[737] = 737;
 buffer[738] = 738;
 buffer[739] = 739;
 buffer[740] = 740;
 buffer[741] = 741;
 buffer[742] = 742;
 buffer[743] = 743;
 buffer[744] = 744;
 buffer[745] = 745;
 buffer[746] = 746;
 buffer[747] = 747;
 buffer[748] = 748;
 buffer[749] = 749;
 buffer[750] = 750;
 buffer[751] = 751;
 buffer[752] = 752;
 buffer[753] = 753;
 buffer[754] = 754;
 buffer[755] = 755;
 buffer[756] = 756;
 buffer[757] = 757;
 buffer[758] = 758;
 buffer[759] = 759;
 buffer[760] = 760;
 buffer[761] = 761;
 buffer[762] = 762;
 buffer[763] = 763;
 buffer[764] = 764;
 buffer[765] = 765;
 buffer[766] = 766;
 buffer[767] = 767;
 buffer[768] = 768;
 buffer[769] = 769;
 buffer[770] = 770;
 buffer[771] = 771;
 buffer[772] = 772;
 buffer[773] = 773;
 buffer[774] = 774;
 buffer[775] = 775;
 buffer[776] = 776;
 buffer[777] = 777;
 buffer[778] = 778;
 buffer[779] = 779;
 buffer[780] = 780;
 buffer[781] = 781;
 buffer[782] = 782;
 buffer[783] = 783;
 buffer[784] = 784;
 buffer[785] = 785;
 buffer[786] = 786;
 buffer[787] = 787;
 buffer[788] = 788;
 buffer[789] = 789;
 buffer[790] = 790;
 buffer[791] = 791;
 buffer[792] = 792;
 buffer[793] = 793;
 buffer[794] = 794;
 buffer[795] = 795;
 buffer[796] = 796;
 buffer[797] = 797;
 buffer[798] = 798;
 buffer[799] = 799;
 buffer[800] = 800;
 buffer[801] = 801;
 buffer[802] = 802;
 buffer[803] = 803;
 buffer[804] = 804;
 buffer[805] = 805;
 buffer[806] = 806;
 buffer[807] = 807;
 buffer[808] = 808;
 buffer[809] = 809;
 buffer[810] = 810;
 buffer[811] = 811;
 buffer[812] = 812;
 buffer[813] = 813;
 buffer[814] = 814;
 buffer[815] = 815;
 buffer[816] = 816;
 buffer[817] = 817;
 buffer[818] = 818;
 buffer[819] = 819;
 buffer[820] = 820;
 buffer[821] = 821;
 buffer[822] = 822;
 buffer[823] = 823;
 buffer[824] = 824;
 buffer[825] = 825;
 buffer[826] = 826;
 buffer[827] = 827;
 buffer[828] = 828;
 buffer[829] = 829;
 buffer[830] = 830;
 buffer[831] = 831;
 buffer[832] = 832;
 buffer[833] = 833;
 buffer[834] = 834;
 buffer[835] = 835;
 buffer[836] = 836;
 buffer[837] = 837;
 buffer[838] = 838;
 buffer[839] = 839;
 buffer[840] = 840;
 buffer[841] = 841;
 buffer[842] = 842;
 buffer[843] = 843;
 buffer[844] = 844;
 buffer[845] = 845;
 buffer[846] = 846;
 buffer[847] = 847;
 buffer[848] = 848;
 buffer[849] = 849;
 buffer[850] = 850;
 buffer[851] = 851;
 buffer[852] = 852;
 buffer[853] = 853;
 buffer[854] = 854;
 buffer[855] = 855;
 buffer[856] = 856;
 buffer[857] = 857;
 buffer[858] = 858;
 buffer[859] = 859;
 buffer[860] = 860;
 buffer[861] = 861;
 buffer[862] = 862;
 buffer[863] = 863;
 buffer[864] = 864;
 buffer[865] = 865;
 buffer[866] = 866;
 buffer[867] = 867;
 buffer[868] = 868;
 buffer[869] = 869;
 buffer[870] = 870;
 buffer[871] = 871;
 buffer[872] = 872;
 buffer[873] = 873;
 buffer[874] = 874;
 buffer[875] = 875;
 buffer[876] = 876;
 buffer[877] = 877;
 buffer[878] = 878;
 buffer[879] = 879;
 buffer[880] = 880;
 buffer[881] = 881;
 buffer[882] = 882;
 buffer[883] = 883;
 buffer[884] = 884;
 buffer[885] = 885;
 buffer[886] = 886;
 buffer[887] = 887;
 buffer[888] = 888;
 buffer[889] = 889;
 buffer[890] = 890;
 buffer[891] = 891;
 buffer[892] = 892;
 buffer[893] = 893;
 buffer[894] = 894;
 buffer[895] = 895;
 buffer[896] = 896;
 buffer[897] = 897;
 buffer[898] = 898;
 buffer[899] = 899;
 buffer[900] = 900;
 buffer[901] = 901;
 buffer[902] = 902;
 buffer[903] = 903;
 buffer[904] = 904;
 buffer[905] = 905;
 buffer[906] = 906;
 buffer[907] = 907;
 buffer[908] = 908;
 buffer[909] = 909;
 buffer[910] = 910;
 buffer[911] = 911;
 buffer[912] = 912;
 buffer[913] = 913;
 buffer[914] = 914;
 buffer[915] = 915;
 buffer[916] = 916;
 buffer[917] = 917;
 buffer[918] = 918;
 buffer[919] = 919;
 buffer[920] = 920;
 buffer[921] = 921;
 buffer[922] = 922;
 buffer[923] = 923;
 buffer[924] = 924;
 buffer[925] = 925;
 buffer[926] = 926;
 buffer[927] = 927;
 buffer[928] = 928;
 buffer[929] = 929;
 buffer[930] = 930;
 buffer[931] = 931;
 buffer[932] = 932;
 buffer[933] = 933;
 buffer[934] = 934;
 buffer[935] = 935;
 buffer[936] = 936;
 buffer[937] = 937;
 buffer[938] = 938;
 buffer[939] = 939;
 buffer[940] = 940;
 buffer[941] = 941;
 buffer[942] = 942;
 buffer[943] = 943;
 buffer[944] = 944;
 buffer[945] = 945;
 buffer[946] = 946;
 buffer[947] = 947;
 buffer[948] = 948;
 buffer[949] = 949;
 buffer[950] = 950;
 buffer[951] = 951;
 buffer[952] = 952;
 buffer[953] = 953;
 buffer[954] = 954;
 buffer[955] = 955;
 buffer[956] = 956;
 buffer[957] = 957;
 buffer[958] = 958;
 buffer[959] = 959;
 buffer[960] = 960;
 buffer[961] = 961;
 buffer[962] = 962;
 buffer[963] = 963;
 buffer[964] = 964;
 buffer[965] = 965;
 buffer[966] = 966;
 buffer[967] = 967;
 buffer[968] = 968;
 buffer[969] = 969;
 buffer[970] = 970;
 buffer[971] = 971;
 buffer[972] = 972;
 buffer[973] = 973;
 buffer[974] = 974;
 buffer[975] = 975;
 buffer[976] = 976;
 buffer[977] = 977;
 buffer[978] = 978;
 buffer[979] = 979;
 buffer[980] = 980;
 buffer[981] = 981;
 buffer[982] = 982;
 buffer[983] = 983;
 buffer[984] = 984;
 buffer[985] = 985;
 buffer[986] = 986;
 buffer[987] = 987;
 buffer[988] = 988;
 buffer[989] = 989;
 buffer[990] = 990;
 buffer[991] = 991;
 buffer[992] = 992;
 buffer[993] = 993;
 buffer[994] = 994;
 buffer[995] = 995;
 buffer[996] = 996;
 buffer[997] = 997;
 buffer[998] = 998;
 buffer[999] = 999;
 buffer[1000] = 1000;
 buffer[1001] = 1001;
 buffer[1002] = 1002;
 buffer[1003] = 1003;
 buffer[1004] = 1004;
 buffer[1005] = 1005;
 buffer[1006] = 1006;
 buffer[1007] = 1007;
 buffer[1008] = 1008;
 buffer[1009] = 1009;
 buffer[1010] = 1010;
 buffer[1011] = 1011;
 buffer[1012] = 1012;
 buffer[1013] = 1013;
 buffer[1014] = 1014;
 buffer[1015] = 1015;
 buffer[1016] = 1016;
 buffer[1017] = 1017;
 buffer[1018] = 1018;
 buffer[1019] = 1019;
 buffer[1020] = 1020;
 buffer[1021] = 1021;
 buffer[1022] = 1022;
 buffer[1023] = 1023;
 buffer[1024] = 1024;
 buffer[1025] = 1025;
 buffer[1026] = 1026;
 buffer[1027] = 1027;
 buffer[1028] = 1028;
 buffer[1029] = 1029;
 buffer[1030] = 1030;
 buffer[1031] = 1031;
 buffer[1032] = 1032;
 buffer[1033] = 1033;
 buffer[1034] = 1034;
 buffer[1035] = 1035;
 buffer[1036] = 1036;
 buffer[1037] = 1037;
 buffer[1038] = 1038;
 buffer[1039] = 1039;
 buffer[1040] = 1040;
 buffer[1041] = 1041;
 buffer[1042] = 1042;
 buffer[1043] = 1043;
 buffer[1044] = 1044;
 buffer[1045] = 1045;
 buffer[1046] = 1046;
 buffer[1047] = 1047;
 buffer[1048] = 1048;
 buffer[1049] = 1049;
 buffer[1050] = 1050;
 buffer[1051] = 1051;
 buffer[1052] = 1052;
 buffer[1053] = 1053;
 buffer[1054] = 1054;
 buffer[1055] = 1055;
 buffer[1056] = 1056;
 buffer[1057] = 1057;
 buffer[1058] = 1058;
 buffer[1059] = 1059;
 buffer[1060] = 1060;
 buffer[1061] = 1061;
 buffer[1062] = 1062;
 buffer[1063] = 1063;
 buffer[1064] = 1064;
 buffer[1065] = 1065;
 buffer[1066] = 1066;
 buffer[1067] = 1067;
 buffer[1068] = 1068;
 buffer[1069] = 1069;
 buffer[1070] = 1070;
 buffer[1071] = 1071;
 buffer[1072] = 1072;
 buffer[1073] = 1073;
 buffer[1074] = 1074;
 buffer[1075] = 1075;
 buffer[1076] = 1076;
 buffer[1077] = 1077;
 buffer[1078] = 1078;
 buffer[1079] = 1079;
 buffer[1080] = 1080;
 buffer[1081] = 1081;
 buffer[1082] = 1082;
 buffer[1083] = 1083;
 buffer[1084] = 1084;
 buffer[1085] = 1085;
 buffer[1086] = 1086;
 buffer[1087] = 1087;
 buffer[1088] = 1088;
 buffer[1089] = 1089;
 buffer[1090] = 1090;
 buffer[1091] = 1091;
 buffer[1092] = 1092;
 buffer[1093] = 1093;
 buffer[1094] = 1094;
 buffer[1095] = 1095;
 buffer[1096] = 1096;
 buffer[1097] = 1097;
 buffer[1098] = 1098;
 buffer[1099] = 1099;
 buffer[1100] = 1100;
 buffer[1101] = 1101;
 buffer[1102] = 1102;
 buffer[1103] = 1103;
 buffer[1104] = 1104;
 buffer[1105] = 1105;
 buffer[1106] = 1106;
 buffer[1107] = 1107;
 buffer[1108] = 1108;
 buffer[1109] = 1109;
 buffer[1110] = 1110;
 buffer[1111] = 1111;
 buffer[1112] = 1112;
 buffer[1113] = 1113;
 buffer[1114] = 1114;
 buffer[1115] = 1115;
 buffer[1116] = 1116;
 buffer[1117] = 1117;
 buffer[1118] = 1118;
 buffer[1119] = 1119;
 buffer[1120] = 1120;
 buffer[1121] = 1121;
 buffer[1122] = 1122;
 buffer[1123] = 1123;
 buffer[1124] = 1124;
 buffer[1125] = 1125;
 buffer[1126] = 1126;
 buffer[1127] = 1127;
 buffer[1128] = 1128;
 buffer[1129] = 1129;
 buffer[1130] = 1130;
 buffer[1131] = 1131;
 buffer[1132] = 1132;
 buffer[1133] = 1133;
 buffer[1134] = 1134;
 buffer[1135] = 1135;
 buffer[1136] = 1136;
 buffer[1137] = 1137;
 buffer[1138] = 1138;
 buffer[1139] = 1139;
 buffer[1140] = 1140;
 buffer[1141] = 1141;
 buffer[1142] = 1142;
 buffer[1143] = 1143;
 buffer[1144] = 1144;
 buffer[1145] = 1145;
 buffer[1146] = 1146;
 buffer[1147] = 1147;
 buffer[1148] = 1148;
 buffer[1149] = 1149;
 buffer[1150] = 1150;
 buffer[1151] = 1151;
 buffer[1152] = 1152;
 buffer[1153] = 1153;
 buffer[1154] = 1154;
 buffer[1155] = 1155;
 buffer[1156] = 1156;
 buffer[1157] = 1157;
 buffer[1158] = 1158;
 buffer[1159] = 1159;
 buffer[1160] = 1160;
 buffer[1161] = 1161;
 buffer[1162] = 1162;
 buffer[1163] = 1163;
 buffer[1164] = 1164;
 buffer[1165] = 1165;
 buffer[1166] = 1166;
 buffer[1167] = 1167;
 buffer[1168] = 1168;
 buffer[1169] = 1169;
 buffer[1170] = 1170;
 buffer[1171] = 1171;
 buffer[1172] = 1172;
 buffer[1173] = 1173;
 buffer[1174] = 1174;
 buffer[1175] = 1175;
 buffer[1176] = 1176;
 buffer[1177] = 1177;
 buffer[1178] = 1178;
 buffer[1179] = 1179;
 buffer[1180] = 1180;
 buffer[1181] = 1181;
 buffer[1182] = 1182;
 buffer[1183] = 1183;
 buffer[1184] = 1184;
 buffer[1185] = 1185;
 buffer[1186] = 1186;
 buffer[1187] = 1187;
 buffer[1188] = 1188;
 buffer[1189] = 1189;
 buffer[1190] = 1190;
 buffer[1191] = 1191;
 buffer[1192] = 1192;
 buffer[1193] = 1193;
 buffer[1194] = 1194;
 buffer[1195] = 1195;
 buffer[1196] = 1196;
 buffer[1197] = 1197;
 buffer[1198] = 1198;
 buffer[1199] = 1199;
 buffer[1200] = 1200;
 buffer[1201] = 1201;
 buffer[1202] = 1202;
 buffer[1203] = 1203;
 buffer[1204] = 1204;
 buffer[1205] = 1205;
 buffer[1206] = 1206;
 buffer[1207] = 1207;
 buffer[1208] = 1208;
 buffer[1209] = 1209;
 buffer[1210] = 1210;
 buffer[1211] = 1211;
 buffer[1212] = 1212;
 buffer[1213] = 1213;
 buffer[1214] = 1214;
 buffer[1215] = 1215;
 buffer[1216] = 1216;
 buffer[1217] = 1217;
 buffer[1218] = 1218;
 buffer[1219] = 1219;
 buffer[1220] = 1220;
 buffer[1221] = 1221;
 buffer[1222] = 1222;
 buffer[1223] = 1223;
 buffer[1224] = 1224;
 buffer[1225] = 1225;
 buffer[1226] = 1226;
 buffer[1227] = 1227;
 buffer[1228] = 1228;
 buffer[1229] = 1229;
 buffer[1230] = 1230;
 buffer[1231] = 1231;
 buffer[1232] = 1232;
 buffer[1233] = 1233;
 buffer[1234] = 1234;
 buffer[1235] = 1235;
 buffer[1236] = 1236;
 buffer[1237] = 1237;
 buffer[1238] = 1238;
 buffer[1239] = 1239;
 buffer[1240] = 1240;
 buffer[1241] = 1241;
 buffer[1242] = 1242;
 buffer[1243] = 1243;
 buffer[1244] = 1244;
 buffer[1245] = 1245;
 buffer[1246] = 1246;
 buffer[1247] = 1247;
 buffer[1248] = 1248;
 buffer[1249] = 1249;
 buffer[1250] = 1250;
 buffer[1251] = 1251;
 buffer[1252] = 1252;
 buffer[1253] = 1253;
 buffer[1254] = 1254;
 buffer[1255] = 1255;
 buffer[1256] = 1256;
 buffer[1257] = 1257;
 buffer[1258] = 1258;
 buffer[1259] = 1259;
 buffer[1260] = 1260;
 buffer[1261] = 1261;
 buffer[1262] = 1262;
 buffer[1263] = 1263;
 buffer[1264] = 1264;
 buffer[1265] = 1265;
 buffer[1266] = 1266;
 buffer[1267] = 1267;
 buffer[1268] = 1268;
 buffer[1269] = 1269;
 buffer[1270] = 1270;
 buffer[1271] = 1271;
 buffer[1272] = 1272;
 buffer[1273] = 1273;
 buffer[1274] = 1274;
 buffer[1275] = 1275;
 buffer[1276] = 1276;
 buffer[1277] = 1277;
 buffer[1278] = 1278;
 buffer[1279] = 1279;
 buffer[1280] = 1280;
 buffer[1281] = 1281;
 buffer[1282] = 1282;
 buffer[1283] = 1283;
 buffer[1284] = 1284;
 buffer[1285] = 1285;
 buffer[1286] = 1286;
 buffer[1287] = 1287;
 buffer[1288] = 1288;
 buffer[1289] = 1289;
 buffer[1290] = 1290;
 buffer[1291] = 1291;
 buffer[1292] = 1292;
 buffer[1293] = 1293;
 buffer[1294] = 1294;
 buffer[1295] = 1295;
 buffer[1296] = 1296;
 buffer[1297] = 1297;
 buffer[1298] = 1298;
 buffer[1299] = 1299;
 buffer[1300] = 1300;
 buffer[1301] = 1301;
 buffer[1302] = 1302;
 buffer[1303] = 1303;
 buffer[1304] = 1304;
 buffer[1305] = 1305;
 buffer[1306] = 1306;
 buffer[1307] = 1307;
 buffer[1308] = 1308;
 buffer[1309] = 1309;
 buffer[1310] = 1310;
 buffer[1311] = 1311;
 buffer[1312] = 1312;
 buffer[1313] = 1313;
 buffer[1314] = 1314;
 buffer[1315] = 1315;
 buffer[1316] = 1316;
 buffer[1317] = 1317;
 buffer[1318] = 1318;
 buffer[1319] = 1319;
 buffer[1320] = 1320;
 buffer[1321] = 1321;
 buffer[1322] = 1322;
 buffer[1323] = 1323;
 buffer[1324] = 1324;
 buffer[1325] = 1325;
 buffer[1326] = 1326;
 buffer[1327] = 1327;
 buffer[1328] = 1328;
 buffer[1329] = 1329;
 buffer[1330] = 1330;
 buffer[1331] = 1331;
 buffer[1332] = 1332;
 buffer[1333] = 1333;
 buffer[1334] = 1334;
 buffer[1335] = 1335;
 buffer[1336] = 1336;
 buffer[1337] = 1337;
 buffer[1338] = 1338;
 buffer[1339] = 1339;
 buffer[1340] = 1340;
 buffer[1341] = 1341;
 buffer[1342] = 1342;
 buffer[1343] = 1343;
 buffer[1344] = 1344;
 buffer[1345] = 1345;
 buffer[1346] = 1346;
 buffer[1347] = 1347;
 buffer[1348] = 1348;
 buffer[1349] = 1349;
 buffer[1350] = 1350;
 buffer[1351] = 1351;
 buffer[1352] = 1352;
 buffer[1353] = 1353;
 buffer[1354] = 1354;
 buffer[1355] = 1355;
 buffer[1356] = 1356;
 buffer[1357] = 1357;
 buffer[1358] = 1358;
 buffer[1359] = 1359;
 buffer[1360] = 1360;
 buffer[1361] = 1361;
 buffer[1362] = 1362;
 buffer[1363] = 1363;
 buffer[1364] = 1364;
 buffer[1365] = 1365;
 buffer[1366] = 1366;
 buffer[1367] = 1367;
 buffer[1368] = 1368;
 buffer[1369] = 1369;
 buffer[1370] = 1370;
 buffer[1371] = 1371;
 buffer[1372] = 1372;
 buffer[1373] = 1373;
 buffer[1374] = 1374;
 buffer[1375] = 1375;
 buffer[1376] = 1376;
 buffer[1377] = 1377;
 buffer[1378] = 1378;
 buffer[1379] = 1379;
 buffer[1380] = 1380;
 buffer[1381] = 1381;
 buffer[1382] = 1382;
 buffer[1383] = 1383;
 buffer[1384] = 1384;
 buffer[1385] = 1385;
 buffer[1386] = 1386;
 buffer[1387] = 1387;
 buffer[1388] = 1388;
 buffer[1389] = 1389;
 buffer[1390] = 1390;
 buffer[1391] = 1391;
 buffer[1392] = 1392;
 buffer[1393] = 1393;
 buffer[1394] = 1394;
 buffer[1395] = 1395;
 buffer[1396] = 1396;
 buffer[1397] = 1397;
 buffer[1398] = 1398;
 buffer[1399] = 1399;
 buffer[1400] = 1400;
 buffer[1401] = 1401;
 buffer[1402] = 1402;
 buffer[1403] = 1403;
 buffer[1404] = 1404;
 buffer[1405] = 1405;
 buffer[1406] = 1406;
 buffer[1407] = 1407;
 buffer[1408] = 1408;
 buffer[1409] = 1409;
 buffer[1410] = 1410;
 buffer[1411] = 1411;
 buffer[1412] = 1412;
 buffer[1413] = 1413;
 buffer[1414] = 1414;
 buffer[1415] = 1415;
 buffer[1416] = 1416;
 buffer[1417] = 1417;
 buffer[1418] = 1418;
 buffer[1419] = 1419;
 buffer[1420] = 1420;
 buffer[1421] = 1421;
 buffer[1422] = 1422;
 buffer[1423] = 1423;
 buffer[1424] = 1424;
 buffer[1425] = 1425;
 buffer[1426] = 1426;
 buffer[1427] = 1427;
 buffer[1428] = 1428;
 buffer[1429] = 1429;
 buffer[1430] = 1430;
 buffer[1431] = 1431;
 buffer[1432] = 1432;
 buffer[1433] = 1433;
 buffer[1434] = 1434;
 buffer[1435] = 1435;
 buffer[1436] = 1436;
 buffer[1437] = 1437;
 buffer[1438] = 1438;
 buffer[1439] = 1439;
 buffer[1440] = 1440;
 buffer[1441] = 1441;
 buffer[1442] = 1442;
 buffer[1443] = 1443;
 buffer[1444] = 1444;
 buffer[1445] = 1445;
 buffer[1446] = 1446;
 buffer[1447] = 1447;
 buffer[1448] = 1448;
 buffer[1449] = 1449;
 buffer[1450] = 1450;
 buffer[1451] = 1451;
 buffer[1452] = 1452;
 buffer[1453] = 1453;
 buffer[1454] = 1454;
 buffer[1455] = 1455;
 buffer[1456] = 1456;
 buffer[1457] = 1457;
 buffer[1458] = 1458;
 buffer[1459] = 1459;
 buffer[1460] = 1460;
 buffer[1461] = 1461;
 buffer[1462] = 1462;
 buffer[1463] = 1463;
 buffer[1464] = 1464;
 buffer[1465] = 1465;
 buffer[1466] = 1466;
 buffer[1467] = 1467;
 buffer[1468] = 1468;
 buffer[1469] = 1469;
 buffer[1470] = 1470;
 buffer[1471] = 1471;
 buffer[1472] = 1472;
 buffer[1473] = 1473;
 buffer[1474] = 1474;
 buffer[1475] = 1475;
 buffer[1476] = 1476;
 buffer[1477] = 1477;
 buffer[1478] = 1478;
 buffer[1479] = 1479;
 buffer[1480] = 1480;
 buffer[1481] = 1481;
 buffer[1482] = 1482;
 buffer[1483] = 1483;
 buffer[1484] = 1484;
 buffer[1485] = 1485;
 buffer[1486] = 1486;
 buffer[1487] = 1487;
 buffer[1488] = 1488;
 buffer[1489] = 1489;
 buffer[1490] = 1490;
 buffer[1491] = 1491;
 buffer[1492] = 1492;
 buffer[1493] = 1493;
 buffer[1494] = 1494;
 buffer[1495] = 1495;
 buffer[1496] = 1496;
 buffer[1497] = 1497;
 buffer[1498] = 1498;
 buffer[1499] = 1499;
 buffer[1500] = 1500;
 buffer[1501] = 1501;
 buffer[1502] = 1502;
 buffer[1503] = 1503;
 buffer[1504] = 1504;
 buffer[1505] = 1505;
 buffer[1506] = 1506;
 buffer[1507] = 1507;
 buffer[1508] = 1508;
 buffer[1509] = 1509;
 buffer[1510] = 1510;
 buffer[1511] = 1511;
 buffer[1512] = 1512;
 buffer[1513] = 1513;
 buffer[1514] = 1514;
 buffer[1515] = 1515;
 buffer[1516] = 1516;
 buffer[1517] = 1517;
 buffer[1518] = 1518;
 buffer[1519] = 1519;
 buffer[1520] = 1520;
 buffer[1521] = 1521;
 buffer[1522] = 1522;
 buffer[1523] = 1523;
 buffer[1524] = 1524;
 buffer[1525] = 1525;
 buffer[1526] = 1526;
 buffer[1527] = 1527;
 buffer[1528] = 1528;
 buffer[1529] = 1529;
 buffer[1530] = 1530;
 buffer[1531] = 1531;
 buffer[1532] = 1532;
 buffer[1533] = 1533;
 buffer[1534] = 1534;
 buffer[1535] = 1535;
 buffer[1536] = 1536;
 buffer[1537] = 1537;
 buffer[1538] = 1538;
 buffer[1539] = 1539;
 buffer[1540] = 1540;
 buffer[1541] = 1541;
 buffer[1542] = 1542;
 buffer[1543] = 1543;
 buffer[1544] = 1544;
 buffer[1545] = 1545;
 buffer[1546] = 1546;
 buffer[1547] = 1547;
 buffer[1548] = 1548;
 buffer[1549] = 1549;
 buffer[1550] = 1550;
 buffer[1551] = 1551;
 buffer[1552] = 1552;
 buffer[1553] = 1553;
 buffer[1554] = 1554;
 buffer[1555] = 1555;
 buffer[1556] = 1556;
 buffer[1557] = 1557;
 buffer[1558] = 1558;
 buffer[1559] = 1559;
 buffer[1560] = 1560;
 buffer[1561] = 1561;
 buffer[1562] = 1562;
 buffer[1563] = 1563;
 buffer[1564] = 1564;
 buffer[1565] = 1565;
 buffer[1566] = 1566;
 buffer[1567] = 1567;
 buffer[1568] = 1568;
 buffer[1569] = 1569;
 buffer[1570] = 1570;
 buffer[1571] = 1571;
 buffer[1572] = 1572;
 buffer[1573] = 1573;
 buffer[1574] = 1574;
 buffer[1575] = 1575;
 buffer[1576] = 1576;
 buffer[1577] = 1577;
 buffer[1578] = 1578;
 buffer[1579] = 1579;
 buffer[1580] = 1580;
 buffer[1581] = 1581;
 buffer[1582] = 1582;
 buffer[1583] = 1583;
 buffer[1584] = 1584;
 buffer[1585] = 1585;
 buffer[1586] = 1586;
 buffer[1587] = 1587;
 buffer[1588] = 1588;
 buffer[1589] = 1589;
 buffer[1590] = 1590;
 buffer[1591] = 1591;
 buffer[1592] = 1592;
 buffer[1593] = 1593;
 buffer[1594] = 1594;
 buffer[1595] = 1595;
 buffer[1596] = 1596;
 buffer[1597] = 1597;
 buffer[1598] = 1598;
 buffer[1599] = 1599;
 buffer[1600] = 1600;
 buffer[1601] = 1601;
 buffer[1602] = 1602;
 buffer[1603] = 1603;
 buffer[1604] = 1604;
 buffer[1605] = 1605;
 buffer[1606] = 1606;
 buffer[1607] = 1607;
 buffer[1608] = 1608;
 buffer[1609] = 1609;
 buffer[1610] = 1610;
 buffer[1611] = 1611;
 buffer[1612] = 1612;
 buffer[1613] = 1613;
 buffer[1614] = 1614;
 buffer[1615] = 1615;
 buffer[1616] = 1616;
 buffer[1617] = 1617;
 buffer[1618] = 1618;
 buffer[1619] = 1619;
 buffer[1620] = 1620;
 buffer[1621] = 1621;
 buffer[1622] = 1622;
 buffer[1623] = 1623;
 buffer[1624] = 1624;
 buffer[1625] = 1625;
 buffer[1626] = 1626;
 buffer[1627] = 1627;
 buffer[1628] = 1628;
 buffer[1629] = 1629;
 buffer[1630] = 1630;
 buffer[1631] = 1631;
 buffer[1632] = 1632;
 buffer[1633] = 1633;
 buffer[1634] = 1634;
 buffer[1635] = 1635;
 buffer[1636] = 1636;
 buffer[1637] = 1637;
 buffer[1638] = 1638;
 buffer[1639] = 1639;
 buffer[1640] = 1640;
 buffer[1641] = 1641;
 buffer[1642] = 1642;
 buffer[1643] = 1643;
 buffer[1644] = 1644;
 buffer[1645] = 1645;
 buffer[1646] = 1646;
 buffer[1647] = 1647;
 buffer[1648] = 1648;
 buffer[1649] = 1649;
 buffer[1650] = 1650;
 buffer[1651] = 1651;
 buffer[1652] = 1652;
 buffer[1653] = 1653;
 buffer[1654] = 1654;
 buffer[1655] = 1655;
 buffer[1656] = 1656;
 buffer[1657] = 1657;
 buffer[1658] = 1658;
 buffer[1659] = 1659;
 buffer[1660] = 1660;
 buffer[1661] = 1661;
 buffer[1662] = 1662;
 buffer[1663] = 1663;
 buffer[1664] = 1664;
 buffer[1665] = 1665;
 buffer[1666] = 1666;
 buffer[1667] = 1667;
 buffer[1668] = 1668;
 buffer[1669] = 1669;
 buffer[1670] = 1670;
 buffer[1671] = 1671;
 buffer[1672] = 1672;
 buffer[1673] = 1673;
 buffer[1674] = 1674;
 buffer[1675] = 1675;
 buffer[1676] = 1676;
 buffer[1677] = 1677;
 buffer[1678] = 1678;
 buffer[1679] = 1679;
 buffer[1680] = 1680;
 buffer[1681] = 1681;
 buffer[1682] = 1682;
 buffer[1683] = 1683;
 buffer[1684] = 1684;
 buffer[1685] = 1685;
 buffer[1686] = 1686;
 buffer[1687] = 1687;
 buffer[1688] = 1688;
 buffer[1689] = 1689;
 buffer[1690] = 1690;
 buffer[1691] = 1691;
 buffer[1692] = 1692;
 buffer[1693] = 1693;
 buffer[1694] = 1694;
 buffer[1695] = 1695;
 buffer[1696] = 1696;
 buffer[1697] = 1697;
 buffer[1698] = 1698;
 buffer[1699] = 1699;
 buffer[1700] = 1700;
 buffer[1701] = 1701;
 buffer[1702] = 1702;
 buffer[1703] = 1703;
 buffer[1704] = 1704;
 buffer[1705] = 1705;
 buffer[1706] = 1706;
 buffer[1707] = 1707;
 buffer[1708] = 1708;
 buffer[1709] = 1709;
 buffer[1710] = 1710;
 buffer[1711] = 1711;
 buffer[1712] = 1712;
 buffer[1713] = 1713;
 buffer[1714] = 1714;
 buffer[1715] = 1715;
 buffer[1716] = 1716;
 buffer[1717] = 1717;
 buffer[1718] = 1718;
 buffer[1719] = 1719;
 buffer[1720] = 1720;
 buffer[1721] = 1721;
 buffer[1722] = 1722;
 buffer[1723] = 1723;
 buffer[1724] = 1724;
 buffer[1725] = 1725;
 buffer[1726] = 1726;
 buffer[1727] = 1727;
 buffer[1728] = 1728;
 buffer[1729] = 1729;
 buffer[1730] = 1730;
 buffer[1731] = 1731;
 buffer[1732] = 1732;
 buffer[1733] = 1733;
 buffer[1734] = 1734;
 buffer[1735] = 1735;
 buffer[1736] = 1736;
 buffer[1737] = 1737;
 buffer[1738] = 1738;
 buffer[1739] = 1739;
 buffer[1740] = 1740;
 buffer[1741] = 1741;
 buffer[1742] = 1742;
 buffer[1743] = 1743;
 buffer[1744] = 1744;
 buffer[1745] = 1745;
 buffer[1746] = 1746;
 buffer[1747] = 1747;
 buffer[1748] = 1748;
 buffer[1749] = 1749;
 buffer[1750] = 1750;
 buffer[1751] = 1751;
 buffer[1752] = 1752;
 buffer[1753] = 1753;
 buffer[1754] = 1754;
 buffer[1755] = 1755;
 buffer[1756] = 1756;
 buffer[1757] = 1757;
 buffer[1758] = 1758;
 buffer[1759] = 1759;
 buffer[1760] = 1760;
 buffer[1761] = 1761;
 buffer[1762] = 1762;
 buffer[1763] = 1763;
 buffer[1764] = 1764;
 buffer[1765] = 1765;
 buffer[1766] = 1766;
 buffer[1767] = 1767;
 buffer[1768] = 1768;
 buffer[1769] = 1769;
 buffer[1770] = 1770;
 buffer[1771] = 1771;
 buffer[1772] = 1772;
 buffer[1773] = 1773;
 buffer[1774] = 1774;
 buffer[1775] = 1775;
 buffer[1776] = 1776;
 buffer[1777] = 1777;
 buffer[1778] = 1778;
 buffer[1779] = 1779;
 buffer[1780] = 1780;
 buffer[1781] = 1781;
 buffer[1782] = 1782;
 buffer[1783] = 1783;
 buffer[1784] = 1784;
 buffer[1785] = 1785;
 buffer[1786] = 1786;
 buffer[1787] = 1787;
 buffer[1788] = 1788;
 buffer[1789] = 1789;
 buffer[1790] = 1790;
 buffer[1791] = 1791;
 buffer[1792] = 1792;
 buffer[1793] = 1793;
 buffer[1794] = 1794;
 buffer[1795] = 1795;
 buffer[1796] = 1796;
 buffer[1797] = 1797;
 buffer[1798] = 1798;
 buffer[1799] = 1799;
 buffer[1800] = 1800;
 buffer[1801] = 1801;
 buffer[1802] = 1802;
 buffer[1803] = 1803;
 buffer[1804] = 1804;
 buffer[1805] = 1805;
 buffer[1806] = 1806;
 buffer[1807] = 1807;
 buffer[1808] = 1808;
 buffer[1809] = 1809;
 buffer[1810] = 1810;
 buffer[1811] = 1811;
 buffer[1812] = 1812;
 buffer[1813] = 1813;
 buffer[1814] = 1814;
 buffer[1815] = 1815;
 buffer[1816] = 1816;
 buffer[1817] = 1817;
 buffer[1818] = 1818;
 buffer[1819] = 1819;
 buffer[1820] = 1820;
 buffer[1821] = 1821;
 buffer[1822] = 1822;
 buffer[1823] = 1823;
 buffer[1824] = 1824;
 buffer[1825] = 1825;
 buffer[1826] = 1826;
 buffer[1827] = 1827;
 buffer[1828] = 1828;
 buffer[1829] = 1829;
 buffer[1830] = 1830;
 buffer[1831] = 1831;
 buffer[1832] = 1832;
 buffer[1833] = 1833;
 buffer[1834] = 1834;
 buffer[1835] = 1835;
 buffer[1836] = 1836;
 buffer[1837] = 1837;
 buffer[1838] = 1838;
 buffer[1839] = 1839;
 buffer[1840] = 1840;
 buffer[1841] = 1841;
 buffer[1842] = 1842;
 buffer[1843] = 1843;
 buffer[1844] = 1844;
 buffer[1845] = 1845;
 buffer[1846] = 1846;
 buffer[1847] = 1847;
 buffer[1848] = 1848;
 buffer[1849] = 1849;
 buffer[1850] = 1850;
 buffer[1851] = 1851;
 buffer[1852] = 1852;
 buffer[1853] = 1853;
 buffer[1854] = 1854;
 buffer[1855] = 1855;
 buffer[1856] = 1856;
 buffer[1857] = 1857;
 buffer[1858] = 1858;
 buffer[1859] = 1859;
 buffer[1860] = 1860;
 buffer[1861] = 1861;
 buffer[1862] = 1862;
 buffer[1863] = 1863;
 buffer[1864] = 1864;
 buffer[1865] = 1865;
 buffer[1866] = 1866;
 buffer[1867] = 1867;
 buffer[1868] = 1868;
 buffer[1869] = 1869;
 buffer[1870] = 1870;
 buffer[1871] = 1871;
 buffer[1872] = 1872;
 buffer[1873] = 1873;
 buffer[1874] = 1874;
 buffer[1875] = 1875;
 buffer[1876] = 1876;
 buffer[1877] = 1877;
 buffer[1878] = 1878;
 buffer[1879] = 1879;
 buffer[1880] = 1880;
 buffer[1881] = 1881;
 buffer[1882] = 1882;
 buffer[1883] = 1883;
 buffer[1884] = 1884;
 buffer[1885] = 1885;
 buffer[1886] = 1886;
 buffer[1887] = 1887;
 buffer[1888] = 1888;
 buffer[1889] = 1889;
 buffer[1890] = 1890;
 buffer[1891] = 1891;
 buffer[1892] = 1892;
 buffer[1893] = 1893;
 buffer[1894] = 1894;
 buffer[1895] = 1895;
 buffer[1896] = 1896;
 buffer[1897] = 1897;
 buffer[1898] = 1898;
 buffer[1899] = 1899;
 buffer[1900] = 1900;
 buffer[1901] = 1901;
 buffer[1902] = 1902;
 buffer[1903] = 1903;
 buffer[1904] = 1904;
 buffer[1905] = 1905;
 buffer[1906] = 1906;
 buffer[1907] = 1907;
 buffer[1908] = 1908;
 buffer[1909] = 1909;
 buffer[1910] = 1910;
 buffer[1911] = 1911;
 buffer[1912] = 1912;
 buffer[1913] = 1913;
 buffer[1914] = 1914;
 buffer[1915] = 1915;
 buffer[1916] = 1916;
 buffer[1917] = 1917;
 buffer[1918] = 1918;
 buffer[1919] = 1919;
 buffer[1920] = 1920;
 buffer[1921] = 1921;
 buffer[1922] = 1922;
 buffer[1923] = 1923;
 buffer[1924] = 1924;
 buffer[1925] = 1925;
 buffer[1926] = 1926;
 buffer[1927] = 1927;
 buffer[1928] = 1928;
 buffer[1929] = 1929;
 buffer[1930] = 1930;
 buffer[1931] = 1931;
 buffer[1932] = 1932;
 buffer[1933] = 1933;
 buffer[1934] = 1934;
 buffer[1935] = 1935;
 buffer[1936] = 1936;
 buffer[1937] = 1937;
 buffer[1938] = 1938;
 buffer[1939] = 1939;
 buffer[1940] = 1940;
 buffer[1941] = 1941;
 buffer[1942] = 1942;
 buffer[1943] = 1943;
 buffer[1944] = 1944;
 buffer[1945] = 1945;
 buffer[1946] = 1946;
 buffer[1947] = 1947;
 buffer[1948] = 1948;
 buffer[1949] = 1949;
 buffer[1950] = 1950;
 buffer[1951] = 1951;
 buffer[1952] = 1952;
 buffer[1953] = 1953;
 buffer[1954] = 1954;
 buffer[1955] = 1955;
 buffer[1956] = 1956;
 buffer[1957] = 1957;
 buffer[1958] = 1958;
 buffer[1959] = 1959;
 buffer[1960] = 1960;
 buffer[1961] = 1961;
 buffer[1962] = 1962;
 buffer[1963] = 1963;
 buffer[1964] = 1964;
 buffer[1965] = 1965;
 buffer[1966] = 1966;
 buffer[1967] = 1967;
 buffer[1968] = 1968;
 buffer[1969] = 1969;
 buffer[1970] = 1970;
 buffer[1971] = 1971;
 buffer[1972] = 1972;
 buffer[1973] = 1973;
 buffer[1974] = 1974;
 buffer[1975] = 1975;
 buffer[1976] = 1976;
 buffer[1977] = 1977;
 buffer[1978] = 1978;
 buffer[1979] = 1979;
 buffer[1980] = 1980;
 buffer[1981] = 1981;
 buffer[1982] = 1982;
 buffer[1983] = 1983;
 buffer[1984] = 1984;
 buffer[1985] = 1985;
 buffer[1986] = 1986;
 buffer[1987] = 1987;
 buffer[1988] = 1988;
 buffer[1989] = 1989;
 buffer[1990] = 1990;
 buffer[1991] = 1991;
 buffer[1992] = 1992;
 buffer[1993] = 1993;
 buffer[1994] = 1994;
 buffer[1995] = 1995;
 buffer[1996] = 1996;
 buffer[1997] = 1997;
 buffer[1998] = 1998;
 buffer[1999] = 1999;
 buffer[2000] = 2000;
 buffer[2001] = 2001;
 buffer[2002] = 2002;
 buffer[2003] = 2003;
 buffer[2004] = 2004;
 buffer[2005] = 2005;
 buffer[2006] = 2006;
 buffer[2007] = 2007;
 buffer[2008] = 2008;
 buffer[2009] = 2009;
 buffer[2010] = 2010;
 buffer[2011] = 2011;
 buffer[2012] = 2012;
 buffer[2013] = 2013;
 buffer[2014] = 2014;
 buffer[2015] = 2015;
 buffer[2016] = 2016;
 buffer[2017] = 2017;
 buffer[2018] = 2018;
 buffer[2019] = 2019;
 buffer[2020] = 2020;
 buffer[2021] = 2021;
 buffer[2022] = 2022;
 buffer[2023] = 2023;
 buffer[2024] = 2024;
 buffer[2025] = 2025;
 buffer[2026] = 2026;
 buffer[2027] = 2027;
 buffer[2028] = 2028;
 buffer[2029] = 2029;
 buffer[2030] = 2030;
 buffer[2031] = 2031;
 buffer[2032] = 2032;
 buffer[2033] = 2033;
 buffer[2034] = 2034;
 buffer[2035] = 2035;
 buffer[2036] = 2036;
 buffer[2037] = 2037;
 buffer[2038] = 2038;
 buffer[2039] = 2039;
 buffer[2040] = 2040;
 buffer[2041] = 2041;
 buffer[2042] = 2042;
 buffer[2043] = 2043;
 buffer[2044] = 2044;
 buffer[2045] = 2045;
 buffer[2046] = 2046;
 buffer[2047] = 2047;
 buffer[2048] = 2048;
 buffer[2049] = 2049;
 buffer[2050] = 2050;
 buffer[2051] = 2051;
 buffer[2052] = 2052;
 buffer[2053] = 2053;
 buffer[2054] = 2054;
 buffer[2055] = 2055;
 buffer[2056] = 2056;
 buffer[2057] = 2057;
 buffer[2058] = 2058;
 buffer[2059] = 2059;
 buffer[2060] = 2060;
 buffer[2061] = 2061;
 buffer[2062] = 2062;
 buffer[2063] = 2063;
 buffer[2064] = 2064;
 buffer[2065] = 2065;
 buffer[2066] = 2066;
 buffer[2067] = 2067;
 buffer[2068] = 2068;
 buffer[2069] = 2069;
 buffer[2070] = 2070;
 buffer[2071] = 2071;
 buffer[2072] = 2072;
 buffer[2073] = 2073;
 buffer[2074] = 2074;
 buffer[2075] = 2075;
 buffer[2076] = 2076;
 buffer[2077] = 2077;
 buffer[2078] = 2078;
 buffer[2079] = 2079;
 buffer[2080] = 2080;
 buffer[2081] = 2081;
 buffer[2082] = 2082;
 buffer[2083] = 2083;
 buffer[2084] = 2084;
 buffer[2085] = 2085;
 buffer[2086] = 2086;
 buffer[2087] = 2087;
 buffer[2088] = 2088;
 buffer[2089] = 2089;
 buffer[2090] = 2090;
 buffer[2091] = 2091;
 buffer[2092] = 2092;
 buffer[2093] = 2093;
 buffer[2094] = 2094;
 buffer[2095] = 2095;
 buffer[2096] = 2096;
 buffer[2097] = 2097;
 buffer[2098] = 2098;
 buffer[2099] = 2099;
 buffer[2100] = 2100;
 buffer[2101] = 2101;
 buffer[2102] = 2102;
 buffer[2103] = 2103;
 buffer[2104] = 2104;
 buffer[2105] = 2105;
 buffer[2106] = 2106;
 buffer[2107] = 2107;
 buffer[2108] = 2108;
 buffer[2109] = 2109;
 buffer[2110] = 2110;
 buffer[2111] = 2111;
 buffer[2112] = 2112;
 buffer[2113] = 2113;
 buffer[2114] = 2114;
 buffer[2115] = 2115;
 buffer[2116] = 2116;
 buffer[2117] = 2117;
 buffer[2118] = 2118;
 buffer[2119] = 2119;
 buffer[2120] = 2120;
 buffer[2121] = 2121;
 buffer[2122] = 2122;
 buffer[2123] = 2123;
 buffer[2124] = 2124;
 buffer[2125] = 2125;
 buffer[2126] = 2126;
 buffer[2127] = 2127;
 buffer[2128] = 2128;
 buffer[2129] = 2129;
 buffer[2130] = 2130;
 buffer[2131] = 2131;
 buffer[2132] = 2132;
 buffer[2133] = 2133;
 buffer[2134] = 2134;
 buffer[2135] = 2135;
 buffer[2136] = 2136;
 buffer[2137] = 2137;
 buffer[2138] = 2138;
 buffer[2139] = 2139;
 buffer[2140] = 2140;
 buffer[2141] = 2141;
 buffer[2142] = 2142;
 buffer[2143] = 2143;
 buffer[2144] = 2144;
 buffer[2145] = 2145;
 buffer[2146] = 2146;
 buffer[2147] = 2147;
 buffer[2148] = 2148;
 buffer[2149] = 2149;
 buffer[2150] = 2150;
 buffer[2151] = 2151;
 buffer[2152] = 2152;
 buffer[2153] = 2153;
 buffer[2154] = 2154;
 buffer[2155] = 2155;
 buffer[2156] = 2156;
 buffer[2157] = 2157;
 buffer[2158] = 2158;
 buffer[2159] = 2159;
 buffer[2160] = 2160;
 buffer[2161] = 2161;
 buffer[2162] = 2162;
 buffer[2163] = 2163;
 buffer[2164] = 2164;
 buffer[2165] = 2165;
 buffer[2166] = 2166;
 buffer[2167] = 2167;
 buffer[2168] = 2168;
 buffer[2169] = 2169;
 buffer[2170] = 2170;
 buffer[2171] = 2171;
 buffer[2172] = 2172;
 buffer[2173] = 2173;
 buffer[2174] = 2174;
 buffer[2175] = 2175;
 buffer[2176] = 2176;
 buffer[2177] = 2177;
 buffer[2178] = 2178;
 buffer[2179] = 2179;
 buffer[2180] = 2180;
 buffer[2181] = 2181;
 buffer[2182] = 2182;
 buffer[2183] = 2183;
 buffer[2184] = 2184;
 buffer[2185] = 2185;
 buffer[2186] = 2186;
 buffer[2187] = 2187;
 buffer[2188] = 2188;
 buffer[2189] = 2189;
 buffer[2190] = 2190;
 buffer[2191] = 2191;
 buffer[2192] = 2192;
 buffer[2193] = 2193;
 buffer[2194] = 2194;
 buffer[2195] = 2195;
 buffer[2196] = 2196;
 buffer[2197] = 2197;
 buffer[2198] = 2198;
 buffer[2199] = 2199;
 buffer[2200] = 2200;
 buffer[2201] = 2201;
 buffer[2202] = 2202;
 buffer[2203] = 2203;
 buffer[2204] = 2204;
 buffer[2205] = 2205;
 buffer[2206] = 2206;
 buffer[2207] = 2207;
 buffer[2208] = 2208;
 buffer[2209] = 2209;
 buffer[2210] = 2210;
 buffer[2211] = 2211;
 buffer[2212] = 2212;
 buffer[2213] = 2213;
 buffer[2214] = 2214;
 buffer[2215] = 2215;
 buffer[2216] = 2216;
 buffer[2217] = 2217;
 buffer[2218] = 2218;
 buffer[2219] = 2219;
 buffer[2220] = 2220;
 buffer[2221] = 2221;
 buffer[2222] = 2222;
 buffer[2223] = 2223;
 buffer[2224] = 2224;
 buffer[2225] = 2225;
 buffer[2226] = 2226;
 buffer[2227] = 2227;
 buffer[2228] = 2228;
 buffer[2229] = 2229;
 buffer[2230] = 2230;
 buffer[2231] = 2231;
 buffer[2232] = 2232;
 buffer[2233] = 2233;
 buffer[2234] = 2234;
 buffer[2235] = 2235;
 buffer[2236] = 2236;
 buffer[2237] = 2237;
 buffer[2238] = 2238;
 buffer[2239] = 2239;
 buffer[2240] = 2240;
 buffer[2241] = 2241;
 buffer[2242] = 2242;
 buffer[2243] = 2243;
 buffer[2244] = 2244;
 buffer[2245] = 2245;
 buffer[2246] = 2246;
 buffer[2247] = 2247;
 buffer[2248] = 2248;
 buffer[2249] = 2249;
 buffer[2250] = 2250;
 buffer[2251] = 2251;
 buffer[2252] = 2252;
 buffer[2253] = 2253;
 buffer[2254] = 2254;
 buffer[2255] = 2255;
 buffer[2256] = 2256;
 buffer[2257] = 2257;
 buffer[2258] = 2258;
 buffer[2259] = 2259;
 buffer[2260] = 2260;
 buffer[2261] = 2261;
 buffer[2262] = 2262;
 buffer[2263] = 2263;
 buffer[2264] = 2264;
 buffer[2265] = 2265;
 buffer[2266] = 2266;
 buffer[2267] = 2267;
 buffer[2268] = 2268;
 buffer[2269] = 2269;
 buffer[2270] = 2270;
 buffer[2271] = 2271;
 buffer[2272] = 2272;
 buffer[2273] = 2273;
 buffer[2274] = 2274;
 buffer[2275] = 2275;
 buffer[2276] = 2276;
 buffer[2277] = 2277;
 buffer[2278] = 2278;
 buffer[2279] = 2279;
 buffer[2280] = 2280;
 buffer[2281] = 2281;
 buffer[2282] = 2282;
 buffer[2283] = 2283;
 buffer[2284] = 2284;
 buffer[2285] = 2285;
 buffer[2286] = 2286;
 buffer[2287] = 2287;
 buffer[2288] = 2288;
 buffer[2289] = 2289;
 buffer[2290] = 2290;
 buffer[2291] = 2291;
 buffer[2292] = 2292;
 buffer[2293] = 2293;
 buffer[2294] = 2294;
 buffer[2295] = 2295;
 buffer[2296] = 2296;
 buffer[2297] = 2297;
 buffer[2298] = 2298;
 buffer[2299] = 2299;
 buffer[2300] = 2300;
 buffer[2301] = 2301;
 buffer[2302] = 2302;
 buffer[2303] = 2303;
 buffer[2304] = 2304;
 buffer[2305] = 2305;
 buffer[2306] = 2306;
 buffer[2307] = 2307;
 buffer[2308] = 2308;
 buffer[2309] = 2309;
 buffer[2310] = 2310;
 buffer[2311] = 2311;
 buffer[2312] = 2312;
 buffer[2313] = 2313;
 buffer[2314] = 2314;
 buffer[2315] = 2315;
 buffer[2316] = 2316;
 buffer[2317] = 2317;
 buffer[2318] = 2318;
 buffer[2319] = 2319;
 buffer[2320] = 2320;
 buffer[2321] = 2321;
 buffer[2322] = 2322;
 buffer[2323] = 2323;
 buffer[2324] = 2324;
 buffer[2325] = 2325;
 buffer[2326] = 2326;
 buffer[2327] = 2327;
 buffer[2328] = 2328;
 buffer[2329] = 2329;
 buffer[2330] = 2330;
 buffer[2331] = 2331;
 buffer[2332] = 2332;
 buffer[2333] = 2333;
 buffer[2334] = 2334;
 buffer[2335] = 2335;
 buffer[2336] = 2336;
 buffer[2337] = 2337;
 buffer[2338] = 2338;
 buffer[2339] = 2339;
 buffer[2340] = 2340;
 buffer[2341] = 2341;
 buffer[2342] = 2342;
 buffer[2343] = 2343;
 buffer[2344] = 2344;
 buffer[2345] = 2345;
 buffer[2346] = 2346;
 buffer[2347] = 2347;
 buffer[2348] = 2348;
 buffer[2349] = 2349;
 buffer[2350] = 2350;
 buffer[2351] = 2351;
 buffer[2352] = 2352;
 buffer[2353] = 2353;
 buffer[2354] = 2354;
 buffer[2355] = 2355;
 buffer[2356] = 2356;
 buffer[2357] = 2357;
 buffer[2358] = 2358;
 buffer[2359] = 2359;
 buffer[2360] = 2360;
 buffer[2361] = 2361;
 buffer[2362] = 2362;
 buffer[2363] = 2363;
 buffer[2364] = 2364;
 buffer[2365] = 2365;
 buffer[2366] = 2366;
 buffer[2367] = 2367;
 buffer[2368] = 2368;
 buffer[2369] = 2369;
 buffer[2370] = 2370;
 buffer[2371] = 2371;
 buffer[2372] = 2372;
 buffer[2373] = 2373;
 buffer[2374] = 2374;
 buffer[2375] = 2375;
 buffer[2376] = 2376;
 buffer[2377] = 2377;
 buffer[2378] = 2378;
 buffer[2379] = 2379;
 buffer[2380] = 2380;
 buffer[2381] = 2381;
 buffer[2382] = 2382;
 buffer[2383] = 2383;
 buffer[2384] = 2384;
 buffer[2385] = 2385;
 buffer[2386] = 2386;
 buffer[2387] = 2387;
 buffer[2388] = 2388;
 buffer[2389] = 2389;
 buffer[2390] = 2390;
 buffer[2391] = 2391;
 buffer[2392] = 2392;
 buffer[2393] = 2393;
 buffer[2394] = 2394;
 buffer[2395] = 2395;
 buffer[2396] = 2396;
 buffer[2397] = 2397;
 buffer[2398] = 2398;
 buffer[2399] = 2399;
end

endmodule

module M_multiplex_display_mem_foreground(
input      [0:0]             in_foreground_wenable0,
input       [7:0]     in_foreground_wdata0,
input      [11:0]                in_foreground_addr0,
input      [0:0]             in_foreground_wenable1,
input      [7:0]                 in_foreground_wdata1,
input      [11:0]                in_foreground_addr1,
output reg  [7:0]     out_foreground_rdata0,
output reg  [7:0]     out_foreground_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2399:0];
always @(posedge clock0) begin
  if (in_foreground_wenable0) begin
    buffer[in_foreground_addr0] <= in_foreground_wdata0;
  end else begin
    out_foreground_rdata0 <= buffer[in_foreground_addr0];
  end
end
always @(posedge clock1) begin
  if (in_foreground_wenable1) begin
    buffer[in_foreground_addr1] <= in_foreground_wdata1;
  end else begin
    out_foreground_rdata1 <= buffer[in_foreground_addr1];
  end
end
initial begin
 buffer[0] = 0;
 buffer[1] = 1;
 buffer[2] = 2;
 buffer[3] = 3;
 buffer[4] = 4;
 buffer[5] = 5;
 buffer[6] = 6;
 buffer[7] = 7;
 buffer[8] = 8;
 buffer[9] = 9;
 buffer[10] = 10;
 buffer[11] = 11;
 buffer[12] = 12;
 buffer[13] = 13;
 buffer[14] = 14;
 buffer[15] = 15;
 buffer[16] = 16;
 buffer[17] = 17;
 buffer[18] = 18;
 buffer[19] = 19;
 buffer[20] = 20;
 buffer[21] = 21;
 buffer[22] = 22;
 buffer[23] = 23;
 buffer[24] = 24;
 buffer[25] = 25;
 buffer[26] = 26;
 buffer[27] = 27;
 buffer[28] = 28;
 buffer[29] = 29;
 buffer[30] = 30;
 buffer[31] = 31;
 buffer[32] = 32;
 buffer[33] = 33;
 buffer[34] = 34;
 buffer[35] = 35;
 buffer[36] = 36;
 buffer[37] = 37;
 buffer[38] = 38;
 buffer[39] = 39;
 buffer[40] = 40;
 buffer[41] = 41;
 buffer[42] = 42;
 buffer[43] = 43;
 buffer[44] = 44;
 buffer[45] = 45;
 buffer[46] = 46;
 buffer[47] = 47;
 buffer[48] = 48;
 buffer[49] = 49;
 buffer[50] = 50;
 buffer[51] = 51;
 buffer[52] = 52;
 buffer[53] = 53;
 buffer[54] = 54;
 buffer[55] = 55;
 buffer[56] = 56;
 buffer[57] = 57;
 buffer[58] = 58;
 buffer[59] = 59;
 buffer[60] = 60;
 buffer[61] = 61;
 buffer[62] = 62;
 buffer[63] = 63;
 buffer[64] = 64;
 buffer[65] = 65;
 buffer[66] = 66;
 buffer[67] = 67;
 buffer[68] = 68;
 buffer[69] = 69;
 buffer[70] = 70;
 buffer[71] = 71;
 buffer[72] = 72;
 buffer[73] = 73;
 buffer[74] = 74;
 buffer[75] = 75;
 buffer[76] = 76;
 buffer[77] = 77;
 buffer[78] = 78;
 buffer[79] = 79;
 buffer[80] = 80;
 buffer[81] = 81;
 buffer[82] = 82;
 buffer[83] = 83;
 buffer[84] = 84;
 buffer[85] = 85;
 buffer[86] = 86;
 buffer[87] = 87;
 buffer[88] = 88;
 buffer[89] = 89;
 buffer[90] = 90;
 buffer[91] = 91;
 buffer[92] = 92;
 buffer[93] = 93;
 buffer[94] = 94;
 buffer[95] = 95;
 buffer[96] = 96;
 buffer[97] = 97;
 buffer[98] = 98;
 buffer[99] = 99;
 buffer[100] = 100;
 buffer[101] = 101;
 buffer[102] = 102;
 buffer[103] = 103;
 buffer[104] = 104;
 buffer[105] = 105;
 buffer[106] = 106;
 buffer[107] = 107;
 buffer[108] = 108;
 buffer[109] = 109;
 buffer[110] = 110;
 buffer[111] = 111;
 buffer[112] = 112;
 buffer[113] = 113;
 buffer[114] = 114;
 buffer[115] = 115;
 buffer[116] = 116;
 buffer[117] = 117;
 buffer[118] = 118;
 buffer[119] = 119;
 buffer[120] = 120;
 buffer[121] = 121;
 buffer[122] = 122;
 buffer[123] = 123;
 buffer[124] = 124;
 buffer[125] = 125;
 buffer[126] = 126;
 buffer[127] = 127;
 buffer[128] = 128;
 buffer[129] = 129;
 buffer[130] = 130;
 buffer[131] = 131;
 buffer[132] = 132;
 buffer[133] = 133;
 buffer[134] = 134;
 buffer[135] = 135;
 buffer[136] = 136;
 buffer[137] = 137;
 buffer[138] = 138;
 buffer[139] = 139;
 buffer[140] = 140;
 buffer[141] = 141;
 buffer[142] = 142;
 buffer[143] = 143;
 buffer[144] = 144;
 buffer[145] = 145;
 buffer[146] = 146;
 buffer[147] = 147;
 buffer[148] = 148;
 buffer[149] = 149;
 buffer[150] = 150;
 buffer[151] = 151;
 buffer[152] = 152;
 buffer[153] = 153;
 buffer[154] = 154;
 buffer[155] = 155;
 buffer[156] = 156;
 buffer[157] = 157;
 buffer[158] = 158;
 buffer[159] = 159;
 buffer[160] = 160;
 buffer[161] = 161;
 buffer[162] = 162;
 buffer[163] = 163;
 buffer[164] = 164;
 buffer[165] = 165;
 buffer[166] = 166;
 buffer[167] = 167;
 buffer[168] = 168;
 buffer[169] = 169;
 buffer[170] = 170;
 buffer[171] = 171;
 buffer[172] = 172;
 buffer[173] = 173;
 buffer[174] = 174;
 buffer[175] = 175;
 buffer[176] = 176;
 buffer[177] = 177;
 buffer[178] = 178;
 buffer[179] = 179;
 buffer[180] = 180;
 buffer[181] = 181;
 buffer[182] = 182;
 buffer[183] = 183;
 buffer[184] = 184;
 buffer[185] = 185;
 buffer[186] = 186;
 buffer[187] = 187;
 buffer[188] = 188;
 buffer[189] = 189;
 buffer[190] = 190;
 buffer[191] = 191;
 buffer[192] = 192;
 buffer[193] = 193;
 buffer[194] = 194;
 buffer[195] = 195;
 buffer[196] = 196;
 buffer[197] = 197;
 buffer[198] = 198;
 buffer[199] = 199;
 buffer[200] = 200;
 buffer[201] = 201;
 buffer[202] = 202;
 buffer[203] = 203;
 buffer[204] = 204;
 buffer[205] = 205;
 buffer[206] = 206;
 buffer[207] = 207;
 buffer[208] = 208;
 buffer[209] = 209;
 buffer[210] = 210;
 buffer[211] = 211;
 buffer[212] = 212;
 buffer[213] = 213;
 buffer[214] = 214;
 buffer[215] = 215;
 buffer[216] = 216;
 buffer[217] = 217;
 buffer[218] = 218;
 buffer[219] = 219;
 buffer[220] = 220;
 buffer[221] = 221;
 buffer[222] = 222;
 buffer[223] = 223;
 buffer[224] = 224;
 buffer[225] = 225;
 buffer[226] = 226;
 buffer[227] = 227;
 buffer[228] = 228;
 buffer[229] = 229;
 buffer[230] = 230;
 buffer[231] = 231;
 buffer[232] = 232;
 buffer[233] = 233;
 buffer[234] = 234;
 buffer[235] = 235;
 buffer[236] = 236;
 buffer[237] = 237;
 buffer[238] = 238;
 buffer[239] = 239;
 buffer[240] = 240;
 buffer[241] = 241;
 buffer[242] = 242;
 buffer[243] = 243;
 buffer[244] = 244;
 buffer[245] = 245;
 buffer[246] = 246;
 buffer[247] = 247;
 buffer[248] = 248;
 buffer[249] = 249;
 buffer[250] = 250;
 buffer[251] = 251;
 buffer[252] = 252;
 buffer[253] = 253;
 buffer[254] = 254;
 buffer[255] = 255;
 buffer[256] = 256;
 buffer[257] = 257;
 buffer[258] = 258;
 buffer[259] = 259;
 buffer[260] = 260;
 buffer[261] = 261;
 buffer[262] = 262;
 buffer[263] = 263;
 buffer[264] = 264;
 buffer[265] = 265;
 buffer[266] = 266;
 buffer[267] = 267;
 buffer[268] = 268;
 buffer[269] = 269;
 buffer[270] = 270;
 buffer[271] = 271;
 buffer[272] = 272;
 buffer[273] = 273;
 buffer[274] = 274;
 buffer[275] = 275;
 buffer[276] = 276;
 buffer[277] = 277;
 buffer[278] = 278;
 buffer[279] = 279;
 buffer[280] = 280;
 buffer[281] = 281;
 buffer[282] = 282;
 buffer[283] = 283;
 buffer[284] = 284;
 buffer[285] = 285;
 buffer[286] = 286;
 buffer[287] = 287;
 buffer[288] = 288;
 buffer[289] = 289;
 buffer[290] = 290;
 buffer[291] = 291;
 buffer[292] = 292;
 buffer[293] = 293;
 buffer[294] = 294;
 buffer[295] = 295;
 buffer[296] = 296;
 buffer[297] = 297;
 buffer[298] = 298;
 buffer[299] = 299;
 buffer[300] = 300;
 buffer[301] = 301;
 buffer[302] = 302;
 buffer[303] = 303;
 buffer[304] = 304;
 buffer[305] = 305;
 buffer[306] = 306;
 buffer[307] = 307;
 buffer[308] = 308;
 buffer[309] = 309;
 buffer[310] = 310;
 buffer[311] = 311;
 buffer[312] = 312;
 buffer[313] = 313;
 buffer[314] = 314;
 buffer[315] = 315;
 buffer[316] = 316;
 buffer[317] = 317;
 buffer[318] = 318;
 buffer[319] = 319;
 buffer[320] = 320;
 buffer[321] = 321;
 buffer[322] = 322;
 buffer[323] = 323;
 buffer[324] = 324;
 buffer[325] = 325;
 buffer[326] = 326;
 buffer[327] = 327;
 buffer[328] = 328;
 buffer[329] = 329;
 buffer[330] = 330;
 buffer[331] = 331;
 buffer[332] = 332;
 buffer[333] = 333;
 buffer[334] = 334;
 buffer[335] = 335;
 buffer[336] = 336;
 buffer[337] = 337;
 buffer[338] = 338;
 buffer[339] = 339;
 buffer[340] = 340;
 buffer[341] = 341;
 buffer[342] = 342;
 buffer[343] = 343;
 buffer[344] = 344;
 buffer[345] = 345;
 buffer[346] = 346;
 buffer[347] = 347;
 buffer[348] = 348;
 buffer[349] = 349;
 buffer[350] = 350;
 buffer[351] = 351;
 buffer[352] = 352;
 buffer[353] = 353;
 buffer[354] = 354;
 buffer[355] = 355;
 buffer[356] = 356;
 buffer[357] = 357;
 buffer[358] = 358;
 buffer[359] = 359;
 buffer[360] = 360;
 buffer[361] = 361;
 buffer[362] = 362;
 buffer[363] = 363;
 buffer[364] = 364;
 buffer[365] = 365;
 buffer[366] = 366;
 buffer[367] = 367;
 buffer[368] = 368;
 buffer[369] = 369;
 buffer[370] = 370;
 buffer[371] = 371;
 buffer[372] = 372;
 buffer[373] = 373;
 buffer[374] = 374;
 buffer[375] = 375;
 buffer[376] = 376;
 buffer[377] = 377;
 buffer[378] = 378;
 buffer[379] = 379;
 buffer[380] = 380;
 buffer[381] = 381;
 buffer[382] = 382;
 buffer[383] = 383;
 buffer[384] = 384;
 buffer[385] = 385;
 buffer[386] = 386;
 buffer[387] = 387;
 buffer[388] = 388;
 buffer[389] = 389;
 buffer[390] = 390;
 buffer[391] = 391;
 buffer[392] = 392;
 buffer[393] = 393;
 buffer[394] = 394;
 buffer[395] = 395;
 buffer[396] = 396;
 buffer[397] = 397;
 buffer[398] = 398;
 buffer[399] = 399;
 buffer[400] = 400;
 buffer[401] = 401;
 buffer[402] = 402;
 buffer[403] = 403;
 buffer[404] = 404;
 buffer[405] = 405;
 buffer[406] = 406;
 buffer[407] = 407;
 buffer[408] = 408;
 buffer[409] = 409;
 buffer[410] = 410;
 buffer[411] = 411;
 buffer[412] = 412;
 buffer[413] = 413;
 buffer[414] = 414;
 buffer[415] = 415;
 buffer[416] = 416;
 buffer[417] = 417;
 buffer[418] = 418;
 buffer[419] = 419;
 buffer[420] = 420;
 buffer[421] = 421;
 buffer[422] = 422;
 buffer[423] = 423;
 buffer[424] = 424;
 buffer[425] = 425;
 buffer[426] = 426;
 buffer[427] = 427;
 buffer[428] = 428;
 buffer[429] = 429;
 buffer[430] = 430;
 buffer[431] = 431;
 buffer[432] = 432;
 buffer[433] = 433;
 buffer[434] = 434;
 buffer[435] = 435;
 buffer[436] = 436;
 buffer[437] = 437;
 buffer[438] = 438;
 buffer[439] = 439;
 buffer[440] = 440;
 buffer[441] = 441;
 buffer[442] = 442;
 buffer[443] = 443;
 buffer[444] = 444;
 buffer[445] = 445;
 buffer[446] = 446;
 buffer[447] = 447;
 buffer[448] = 448;
 buffer[449] = 449;
 buffer[450] = 450;
 buffer[451] = 451;
 buffer[452] = 452;
 buffer[453] = 453;
 buffer[454] = 454;
 buffer[455] = 455;
 buffer[456] = 456;
 buffer[457] = 457;
 buffer[458] = 458;
 buffer[459] = 459;
 buffer[460] = 460;
 buffer[461] = 461;
 buffer[462] = 462;
 buffer[463] = 463;
 buffer[464] = 464;
 buffer[465] = 465;
 buffer[466] = 466;
 buffer[467] = 467;
 buffer[468] = 468;
 buffer[469] = 469;
 buffer[470] = 470;
 buffer[471] = 471;
 buffer[472] = 472;
 buffer[473] = 473;
 buffer[474] = 474;
 buffer[475] = 475;
 buffer[476] = 476;
 buffer[477] = 477;
 buffer[478] = 478;
 buffer[479] = 479;
 buffer[480] = 480;
 buffer[481] = 481;
 buffer[482] = 482;
 buffer[483] = 483;
 buffer[484] = 484;
 buffer[485] = 485;
 buffer[486] = 486;
 buffer[487] = 487;
 buffer[488] = 488;
 buffer[489] = 489;
 buffer[490] = 490;
 buffer[491] = 491;
 buffer[492] = 492;
 buffer[493] = 493;
 buffer[494] = 494;
 buffer[495] = 495;
 buffer[496] = 496;
 buffer[497] = 497;
 buffer[498] = 498;
 buffer[499] = 499;
 buffer[500] = 500;
 buffer[501] = 501;
 buffer[502] = 502;
 buffer[503] = 503;
 buffer[504] = 504;
 buffer[505] = 505;
 buffer[506] = 506;
 buffer[507] = 507;
 buffer[508] = 508;
 buffer[509] = 509;
 buffer[510] = 510;
 buffer[511] = 511;
 buffer[512] = 512;
 buffer[513] = 513;
 buffer[514] = 514;
 buffer[515] = 515;
 buffer[516] = 516;
 buffer[517] = 517;
 buffer[518] = 518;
 buffer[519] = 519;
 buffer[520] = 520;
 buffer[521] = 521;
 buffer[522] = 522;
 buffer[523] = 523;
 buffer[524] = 524;
 buffer[525] = 525;
 buffer[526] = 526;
 buffer[527] = 527;
 buffer[528] = 528;
 buffer[529] = 529;
 buffer[530] = 530;
 buffer[531] = 531;
 buffer[532] = 532;
 buffer[533] = 533;
 buffer[534] = 534;
 buffer[535] = 535;
 buffer[536] = 536;
 buffer[537] = 537;
 buffer[538] = 538;
 buffer[539] = 539;
 buffer[540] = 540;
 buffer[541] = 541;
 buffer[542] = 542;
 buffer[543] = 543;
 buffer[544] = 544;
 buffer[545] = 545;
 buffer[546] = 546;
 buffer[547] = 547;
 buffer[548] = 548;
 buffer[549] = 549;
 buffer[550] = 550;
 buffer[551] = 551;
 buffer[552] = 552;
 buffer[553] = 553;
 buffer[554] = 554;
 buffer[555] = 555;
 buffer[556] = 556;
 buffer[557] = 557;
 buffer[558] = 558;
 buffer[559] = 559;
 buffer[560] = 560;
 buffer[561] = 561;
 buffer[562] = 562;
 buffer[563] = 563;
 buffer[564] = 564;
 buffer[565] = 565;
 buffer[566] = 566;
 buffer[567] = 567;
 buffer[568] = 568;
 buffer[569] = 569;
 buffer[570] = 570;
 buffer[571] = 571;
 buffer[572] = 572;
 buffer[573] = 573;
 buffer[574] = 574;
 buffer[575] = 575;
 buffer[576] = 576;
 buffer[577] = 577;
 buffer[578] = 578;
 buffer[579] = 579;
 buffer[580] = 580;
 buffer[581] = 581;
 buffer[582] = 582;
 buffer[583] = 583;
 buffer[584] = 584;
 buffer[585] = 585;
 buffer[586] = 586;
 buffer[587] = 587;
 buffer[588] = 588;
 buffer[589] = 589;
 buffer[590] = 590;
 buffer[591] = 591;
 buffer[592] = 592;
 buffer[593] = 593;
 buffer[594] = 594;
 buffer[595] = 595;
 buffer[596] = 596;
 buffer[597] = 597;
 buffer[598] = 598;
 buffer[599] = 599;
 buffer[600] = 600;
 buffer[601] = 601;
 buffer[602] = 602;
 buffer[603] = 603;
 buffer[604] = 604;
 buffer[605] = 605;
 buffer[606] = 606;
 buffer[607] = 607;
 buffer[608] = 608;
 buffer[609] = 609;
 buffer[610] = 610;
 buffer[611] = 611;
 buffer[612] = 612;
 buffer[613] = 613;
 buffer[614] = 614;
 buffer[615] = 615;
 buffer[616] = 616;
 buffer[617] = 617;
 buffer[618] = 618;
 buffer[619] = 619;
 buffer[620] = 620;
 buffer[621] = 621;
 buffer[622] = 622;
 buffer[623] = 623;
 buffer[624] = 624;
 buffer[625] = 625;
 buffer[626] = 626;
 buffer[627] = 627;
 buffer[628] = 628;
 buffer[629] = 629;
 buffer[630] = 630;
 buffer[631] = 631;
 buffer[632] = 632;
 buffer[633] = 633;
 buffer[634] = 634;
 buffer[635] = 635;
 buffer[636] = 636;
 buffer[637] = 637;
 buffer[638] = 638;
 buffer[639] = 639;
 buffer[640] = 640;
 buffer[641] = 641;
 buffer[642] = 642;
 buffer[643] = 643;
 buffer[644] = 644;
 buffer[645] = 645;
 buffer[646] = 646;
 buffer[647] = 647;
 buffer[648] = 648;
 buffer[649] = 649;
 buffer[650] = 650;
 buffer[651] = 651;
 buffer[652] = 652;
 buffer[653] = 653;
 buffer[654] = 654;
 buffer[655] = 655;
 buffer[656] = 656;
 buffer[657] = 657;
 buffer[658] = 658;
 buffer[659] = 659;
 buffer[660] = 660;
 buffer[661] = 661;
 buffer[662] = 662;
 buffer[663] = 663;
 buffer[664] = 664;
 buffer[665] = 665;
 buffer[666] = 666;
 buffer[667] = 667;
 buffer[668] = 668;
 buffer[669] = 669;
 buffer[670] = 670;
 buffer[671] = 671;
 buffer[672] = 672;
 buffer[673] = 673;
 buffer[674] = 674;
 buffer[675] = 675;
 buffer[676] = 676;
 buffer[677] = 677;
 buffer[678] = 678;
 buffer[679] = 679;
 buffer[680] = 680;
 buffer[681] = 681;
 buffer[682] = 682;
 buffer[683] = 683;
 buffer[684] = 684;
 buffer[685] = 685;
 buffer[686] = 686;
 buffer[687] = 687;
 buffer[688] = 688;
 buffer[689] = 689;
 buffer[690] = 690;
 buffer[691] = 691;
 buffer[692] = 692;
 buffer[693] = 693;
 buffer[694] = 694;
 buffer[695] = 695;
 buffer[696] = 696;
 buffer[697] = 697;
 buffer[698] = 698;
 buffer[699] = 699;
 buffer[700] = 700;
 buffer[701] = 701;
 buffer[702] = 702;
 buffer[703] = 703;
 buffer[704] = 704;
 buffer[705] = 705;
 buffer[706] = 706;
 buffer[707] = 707;
 buffer[708] = 708;
 buffer[709] = 709;
 buffer[710] = 710;
 buffer[711] = 711;
 buffer[712] = 712;
 buffer[713] = 713;
 buffer[714] = 714;
 buffer[715] = 715;
 buffer[716] = 716;
 buffer[717] = 717;
 buffer[718] = 718;
 buffer[719] = 719;
 buffer[720] = 720;
 buffer[721] = 721;
 buffer[722] = 722;
 buffer[723] = 723;
 buffer[724] = 724;
 buffer[725] = 725;
 buffer[726] = 726;
 buffer[727] = 727;
 buffer[728] = 728;
 buffer[729] = 729;
 buffer[730] = 730;
 buffer[731] = 731;
 buffer[732] = 732;
 buffer[733] = 733;
 buffer[734] = 734;
 buffer[735] = 735;
 buffer[736] = 736;
 buffer[737] = 737;
 buffer[738] = 738;
 buffer[739] = 739;
 buffer[740] = 740;
 buffer[741] = 741;
 buffer[742] = 742;
 buffer[743] = 743;
 buffer[744] = 744;
 buffer[745] = 745;
 buffer[746] = 746;
 buffer[747] = 747;
 buffer[748] = 748;
 buffer[749] = 749;
 buffer[750] = 750;
 buffer[751] = 751;
 buffer[752] = 752;
 buffer[753] = 753;
 buffer[754] = 754;
 buffer[755] = 755;
 buffer[756] = 756;
 buffer[757] = 757;
 buffer[758] = 758;
 buffer[759] = 759;
 buffer[760] = 760;
 buffer[761] = 761;
 buffer[762] = 762;
 buffer[763] = 763;
 buffer[764] = 764;
 buffer[765] = 765;
 buffer[766] = 766;
 buffer[767] = 767;
 buffer[768] = 768;
 buffer[769] = 769;
 buffer[770] = 770;
 buffer[771] = 771;
 buffer[772] = 772;
 buffer[773] = 773;
 buffer[774] = 774;
 buffer[775] = 775;
 buffer[776] = 776;
 buffer[777] = 777;
 buffer[778] = 778;
 buffer[779] = 779;
 buffer[780] = 780;
 buffer[781] = 781;
 buffer[782] = 782;
 buffer[783] = 783;
 buffer[784] = 784;
 buffer[785] = 785;
 buffer[786] = 786;
 buffer[787] = 787;
 buffer[788] = 788;
 buffer[789] = 789;
 buffer[790] = 790;
 buffer[791] = 791;
 buffer[792] = 792;
 buffer[793] = 793;
 buffer[794] = 794;
 buffer[795] = 795;
 buffer[796] = 796;
 buffer[797] = 797;
 buffer[798] = 798;
 buffer[799] = 799;
 buffer[800] = 800;
 buffer[801] = 801;
 buffer[802] = 802;
 buffer[803] = 803;
 buffer[804] = 804;
 buffer[805] = 805;
 buffer[806] = 806;
 buffer[807] = 807;
 buffer[808] = 808;
 buffer[809] = 809;
 buffer[810] = 810;
 buffer[811] = 811;
 buffer[812] = 812;
 buffer[813] = 813;
 buffer[814] = 814;
 buffer[815] = 815;
 buffer[816] = 816;
 buffer[817] = 817;
 buffer[818] = 818;
 buffer[819] = 819;
 buffer[820] = 820;
 buffer[821] = 821;
 buffer[822] = 822;
 buffer[823] = 823;
 buffer[824] = 824;
 buffer[825] = 825;
 buffer[826] = 826;
 buffer[827] = 827;
 buffer[828] = 828;
 buffer[829] = 829;
 buffer[830] = 830;
 buffer[831] = 831;
 buffer[832] = 832;
 buffer[833] = 833;
 buffer[834] = 834;
 buffer[835] = 835;
 buffer[836] = 836;
 buffer[837] = 837;
 buffer[838] = 838;
 buffer[839] = 839;
 buffer[840] = 840;
 buffer[841] = 841;
 buffer[842] = 842;
 buffer[843] = 843;
 buffer[844] = 844;
 buffer[845] = 845;
 buffer[846] = 846;
 buffer[847] = 847;
 buffer[848] = 848;
 buffer[849] = 849;
 buffer[850] = 850;
 buffer[851] = 851;
 buffer[852] = 852;
 buffer[853] = 853;
 buffer[854] = 854;
 buffer[855] = 855;
 buffer[856] = 856;
 buffer[857] = 857;
 buffer[858] = 858;
 buffer[859] = 859;
 buffer[860] = 860;
 buffer[861] = 861;
 buffer[862] = 862;
 buffer[863] = 863;
 buffer[864] = 864;
 buffer[865] = 865;
 buffer[866] = 866;
 buffer[867] = 867;
 buffer[868] = 868;
 buffer[869] = 869;
 buffer[870] = 870;
 buffer[871] = 871;
 buffer[872] = 872;
 buffer[873] = 873;
 buffer[874] = 874;
 buffer[875] = 875;
 buffer[876] = 876;
 buffer[877] = 877;
 buffer[878] = 878;
 buffer[879] = 879;
 buffer[880] = 880;
 buffer[881] = 881;
 buffer[882] = 882;
 buffer[883] = 883;
 buffer[884] = 884;
 buffer[885] = 885;
 buffer[886] = 886;
 buffer[887] = 887;
 buffer[888] = 888;
 buffer[889] = 889;
 buffer[890] = 890;
 buffer[891] = 891;
 buffer[892] = 892;
 buffer[893] = 893;
 buffer[894] = 894;
 buffer[895] = 895;
 buffer[896] = 896;
 buffer[897] = 897;
 buffer[898] = 898;
 buffer[899] = 899;
 buffer[900] = 900;
 buffer[901] = 901;
 buffer[902] = 902;
 buffer[903] = 903;
 buffer[904] = 904;
 buffer[905] = 905;
 buffer[906] = 906;
 buffer[907] = 907;
 buffer[908] = 908;
 buffer[909] = 909;
 buffer[910] = 910;
 buffer[911] = 911;
 buffer[912] = 912;
 buffer[913] = 913;
 buffer[914] = 914;
 buffer[915] = 915;
 buffer[916] = 916;
 buffer[917] = 917;
 buffer[918] = 918;
 buffer[919] = 919;
 buffer[920] = 920;
 buffer[921] = 921;
 buffer[922] = 922;
 buffer[923] = 923;
 buffer[924] = 924;
 buffer[925] = 925;
 buffer[926] = 926;
 buffer[927] = 927;
 buffer[928] = 928;
 buffer[929] = 929;
 buffer[930] = 930;
 buffer[931] = 931;
 buffer[932] = 932;
 buffer[933] = 933;
 buffer[934] = 934;
 buffer[935] = 935;
 buffer[936] = 936;
 buffer[937] = 937;
 buffer[938] = 938;
 buffer[939] = 939;
 buffer[940] = 940;
 buffer[941] = 941;
 buffer[942] = 942;
 buffer[943] = 943;
 buffer[944] = 944;
 buffer[945] = 945;
 buffer[946] = 946;
 buffer[947] = 947;
 buffer[948] = 948;
 buffer[949] = 949;
 buffer[950] = 950;
 buffer[951] = 951;
 buffer[952] = 952;
 buffer[953] = 953;
 buffer[954] = 954;
 buffer[955] = 955;
 buffer[956] = 956;
 buffer[957] = 957;
 buffer[958] = 958;
 buffer[959] = 959;
 buffer[960] = 960;
 buffer[961] = 961;
 buffer[962] = 962;
 buffer[963] = 963;
 buffer[964] = 964;
 buffer[965] = 965;
 buffer[966] = 966;
 buffer[967] = 967;
 buffer[968] = 968;
 buffer[969] = 969;
 buffer[970] = 970;
 buffer[971] = 971;
 buffer[972] = 972;
 buffer[973] = 973;
 buffer[974] = 974;
 buffer[975] = 975;
 buffer[976] = 976;
 buffer[977] = 977;
 buffer[978] = 978;
 buffer[979] = 979;
 buffer[980] = 980;
 buffer[981] = 981;
 buffer[982] = 982;
 buffer[983] = 983;
 buffer[984] = 984;
 buffer[985] = 985;
 buffer[986] = 986;
 buffer[987] = 987;
 buffer[988] = 988;
 buffer[989] = 989;
 buffer[990] = 990;
 buffer[991] = 991;
 buffer[992] = 992;
 buffer[993] = 993;
 buffer[994] = 994;
 buffer[995] = 995;
 buffer[996] = 996;
 buffer[997] = 997;
 buffer[998] = 998;
 buffer[999] = 999;
 buffer[1000] = 1000;
 buffer[1001] = 1001;
 buffer[1002] = 1002;
 buffer[1003] = 1003;
 buffer[1004] = 1004;
 buffer[1005] = 1005;
 buffer[1006] = 1006;
 buffer[1007] = 1007;
 buffer[1008] = 1008;
 buffer[1009] = 1009;
 buffer[1010] = 1010;
 buffer[1011] = 1011;
 buffer[1012] = 1012;
 buffer[1013] = 1013;
 buffer[1014] = 1014;
 buffer[1015] = 1015;
 buffer[1016] = 1016;
 buffer[1017] = 1017;
 buffer[1018] = 1018;
 buffer[1019] = 1019;
 buffer[1020] = 1020;
 buffer[1021] = 1021;
 buffer[1022] = 1022;
 buffer[1023] = 1023;
 buffer[1024] = 1024;
 buffer[1025] = 1025;
 buffer[1026] = 1026;
 buffer[1027] = 1027;
 buffer[1028] = 1028;
 buffer[1029] = 1029;
 buffer[1030] = 1030;
 buffer[1031] = 1031;
 buffer[1032] = 1032;
 buffer[1033] = 1033;
 buffer[1034] = 1034;
 buffer[1035] = 1035;
 buffer[1036] = 1036;
 buffer[1037] = 1037;
 buffer[1038] = 1038;
 buffer[1039] = 1039;
 buffer[1040] = 1040;
 buffer[1041] = 1041;
 buffer[1042] = 1042;
 buffer[1043] = 1043;
 buffer[1044] = 1044;
 buffer[1045] = 1045;
 buffer[1046] = 1046;
 buffer[1047] = 1047;
 buffer[1048] = 1048;
 buffer[1049] = 1049;
 buffer[1050] = 1050;
 buffer[1051] = 1051;
 buffer[1052] = 1052;
 buffer[1053] = 1053;
 buffer[1054] = 1054;
 buffer[1055] = 1055;
 buffer[1056] = 1056;
 buffer[1057] = 1057;
 buffer[1058] = 1058;
 buffer[1059] = 1059;
 buffer[1060] = 1060;
 buffer[1061] = 1061;
 buffer[1062] = 1062;
 buffer[1063] = 1063;
 buffer[1064] = 1064;
 buffer[1065] = 1065;
 buffer[1066] = 1066;
 buffer[1067] = 1067;
 buffer[1068] = 1068;
 buffer[1069] = 1069;
 buffer[1070] = 1070;
 buffer[1071] = 1071;
 buffer[1072] = 1072;
 buffer[1073] = 1073;
 buffer[1074] = 1074;
 buffer[1075] = 1075;
 buffer[1076] = 1076;
 buffer[1077] = 1077;
 buffer[1078] = 1078;
 buffer[1079] = 1079;
 buffer[1080] = 1080;
 buffer[1081] = 1081;
 buffer[1082] = 1082;
 buffer[1083] = 1083;
 buffer[1084] = 1084;
 buffer[1085] = 1085;
 buffer[1086] = 1086;
 buffer[1087] = 1087;
 buffer[1088] = 1088;
 buffer[1089] = 1089;
 buffer[1090] = 1090;
 buffer[1091] = 1091;
 buffer[1092] = 1092;
 buffer[1093] = 1093;
 buffer[1094] = 1094;
 buffer[1095] = 1095;
 buffer[1096] = 1096;
 buffer[1097] = 1097;
 buffer[1098] = 1098;
 buffer[1099] = 1099;
 buffer[1100] = 1100;
 buffer[1101] = 1101;
 buffer[1102] = 1102;
 buffer[1103] = 1103;
 buffer[1104] = 1104;
 buffer[1105] = 1105;
 buffer[1106] = 1106;
 buffer[1107] = 1107;
 buffer[1108] = 1108;
 buffer[1109] = 1109;
 buffer[1110] = 1110;
 buffer[1111] = 1111;
 buffer[1112] = 1112;
 buffer[1113] = 1113;
 buffer[1114] = 1114;
 buffer[1115] = 1115;
 buffer[1116] = 1116;
 buffer[1117] = 1117;
 buffer[1118] = 1118;
 buffer[1119] = 1119;
 buffer[1120] = 1120;
 buffer[1121] = 1121;
 buffer[1122] = 1122;
 buffer[1123] = 1123;
 buffer[1124] = 1124;
 buffer[1125] = 1125;
 buffer[1126] = 1126;
 buffer[1127] = 1127;
 buffer[1128] = 1128;
 buffer[1129] = 1129;
 buffer[1130] = 1130;
 buffer[1131] = 1131;
 buffer[1132] = 1132;
 buffer[1133] = 1133;
 buffer[1134] = 1134;
 buffer[1135] = 1135;
 buffer[1136] = 1136;
 buffer[1137] = 1137;
 buffer[1138] = 1138;
 buffer[1139] = 1139;
 buffer[1140] = 1140;
 buffer[1141] = 1141;
 buffer[1142] = 1142;
 buffer[1143] = 1143;
 buffer[1144] = 1144;
 buffer[1145] = 1145;
 buffer[1146] = 1146;
 buffer[1147] = 1147;
 buffer[1148] = 1148;
 buffer[1149] = 1149;
 buffer[1150] = 1150;
 buffer[1151] = 1151;
 buffer[1152] = 1152;
 buffer[1153] = 1153;
 buffer[1154] = 1154;
 buffer[1155] = 1155;
 buffer[1156] = 1156;
 buffer[1157] = 1157;
 buffer[1158] = 1158;
 buffer[1159] = 1159;
 buffer[1160] = 1160;
 buffer[1161] = 1161;
 buffer[1162] = 1162;
 buffer[1163] = 1163;
 buffer[1164] = 1164;
 buffer[1165] = 1165;
 buffer[1166] = 1166;
 buffer[1167] = 1167;
 buffer[1168] = 1168;
 buffer[1169] = 1169;
 buffer[1170] = 1170;
 buffer[1171] = 1171;
 buffer[1172] = 1172;
 buffer[1173] = 1173;
 buffer[1174] = 1174;
 buffer[1175] = 1175;
 buffer[1176] = 1176;
 buffer[1177] = 1177;
 buffer[1178] = 1178;
 buffer[1179] = 1179;
 buffer[1180] = 1180;
 buffer[1181] = 1181;
 buffer[1182] = 1182;
 buffer[1183] = 1183;
 buffer[1184] = 1184;
 buffer[1185] = 1185;
 buffer[1186] = 1186;
 buffer[1187] = 1187;
 buffer[1188] = 1188;
 buffer[1189] = 1189;
 buffer[1190] = 1190;
 buffer[1191] = 1191;
 buffer[1192] = 1192;
 buffer[1193] = 1193;
 buffer[1194] = 1194;
 buffer[1195] = 1195;
 buffer[1196] = 1196;
 buffer[1197] = 1197;
 buffer[1198] = 1198;
 buffer[1199] = 1199;
 buffer[1200] = 1200;
 buffer[1201] = 1201;
 buffer[1202] = 1202;
 buffer[1203] = 1203;
 buffer[1204] = 1204;
 buffer[1205] = 1205;
 buffer[1206] = 1206;
 buffer[1207] = 1207;
 buffer[1208] = 1208;
 buffer[1209] = 1209;
 buffer[1210] = 1210;
 buffer[1211] = 1211;
 buffer[1212] = 1212;
 buffer[1213] = 1213;
 buffer[1214] = 1214;
 buffer[1215] = 1215;
 buffer[1216] = 1216;
 buffer[1217] = 1217;
 buffer[1218] = 1218;
 buffer[1219] = 1219;
 buffer[1220] = 1220;
 buffer[1221] = 1221;
 buffer[1222] = 1222;
 buffer[1223] = 1223;
 buffer[1224] = 1224;
 buffer[1225] = 1225;
 buffer[1226] = 1226;
 buffer[1227] = 1227;
 buffer[1228] = 1228;
 buffer[1229] = 1229;
 buffer[1230] = 1230;
 buffer[1231] = 1231;
 buffer[1232] = 1232;
 buffer[1233] = 1233;
 buffer[1234] = 1234;
 buffer[1235] = 1235;
 buffer[1236] = 1236;
 buffer[1237] = 1237;
 buffer[1238] = 1238;
 buffer[1239] = 1239;
 buffer[1240] = 1240;
 buffer[1241] = 1241;
 buffer[1242] = 1242;
 buffer[1243] = 1243;
 buffer[1244] = 1244;
 buffer[1245] = 1245;
 buffer[1246] = 1246;
 buffer[1247] = 1247;
 buffer[1248] = 1248;
 buffer[1249] = 1249;
 buffer[1250] = 1250;
 buffer[1251] = 1251;
 buffer[1252] = 1252;
 buffer[1253] = 1253;
 buffer[1254] = 1254;
 buffer[1255] = 1255;
 buffer[1256] = 1256;
 buffer[1257] = 1257;
 buffer[1258] = 1258;
 buffer[1259] = 1259;
 buffer[1260] = 1260;
 buffer[1261] = 1261;
 buffer[1262] = 1262;
 buffer[1263] = 1263;
 buffer[1264] = 1264;
 buffer[1265] = 1265;
 buffer[1266] = 1266;
 buffer[1267] = 1267;
 buffer[1268] = 1268;
 buffer[1269] = 1269;
 buffer[1270] = 1270;
 buffer[1271] = 1271;
 buffer[1272] = 1272;
 buffer[1273] = 1273;
 buffer[1274] = 1274;
 buffer[1275] = 1275;
 buffer[1276] = 1276;
 buffer[1277] = 1277;
 buffer[1278] = 1278;
 buffer[1279] = 1279;
 buffer[1280] = 1280;
 buffer[1281] = 1281;
 buffer[1282] = 1282;
 buffer[1283] = 1283;
 buffer[1284] = 1284;
 buffer[1285] = 1285;
 buffer[1286] = 1286;
 buffer[1287] = 1287;
 buffer[1288] = 1288;
 buffer[1289] = 1289;
 buffer[1290] = 1290;
 buffer[1291] = 1291;
 buffer[1292] = 1292;
 buffer[1293] = 1293;
 buffer[1294] = 1294;
 buffer[1295] = 1295;
 buffer[1296] = 1296;
 buffer[1297] = 1297;
 buffer[1298] = 1298;
 buffer[1299] = 1299;
 buffer[1300] = 1300;
 buffer[1301] = 1301;
 buffer[1302] = 1302;
 buffer[1303] = 1303;
 buffer[1304] = 1304;
 buffer[1305] = 1305;
 buffer[1306] = 1306;
 buffer[1307] = 1307;
 buffer[1308] = 1308;
 buffer[1309] = 1309;
 buffer[1310] = 1310;
 buffer[1311] = 1311;
 buffer[1312] = 1312;
 buffer[1313] = 1313;
 buffer[1314] = 1314;
 buffer[1315] = 1315;
 buffer[1316] = 1316;
 buffer[1317] = 1317;
 buffer[1318] = 1318;
 buffer[1319] = 1319;
 buffer[1320] = 1320;
 buffer[1321] = 1321;
 buffer[1322] = 1322;
 buffer[1323] = 1323;
 buffer[1324] = 1324;
 buffer[1325] = 1325;
 buffer[1326] = 1326;
 buffer[1327] = 1327;
 buffer[1328] = 1328;
 buffer[1329] = 1329;
 buffer[1330] = 1330;
 buffer[1331] = 1331;
 buffer[1332] = 1332;
 buffer[1333] = 1333;
 buffer[1334] = 1334;
 buffer[1335] = 1335;
 buffer[1336] = 1336;
 buffer[1337] = 1337;
 buffer[1338] = 1338;
 buffer[1339] = 1339;
 buffer[1340] = 1340;
 buffer[1341] = 1341;
 buffer[1342] = 1342;
 buffer[1343] = 1343;
 buffer[1344] = 1344;
 buffer[1345] = 1345;
 buffer[1346] = 1346;
 buffer[1347] = 1347;
 buffer[1348] = 1348;
 buffer[1349] = 1349;
 buffer[1350] = 1350;
 buffer[1351] = 1351;
 buffer[1352] = 1352;
 buffer[1353] = 1353;
 buffer[1354] = 1354;
 buffer[1355] = 1355;
 buffer[1356] = 1356;
 buffer[1357] = 1357;
 buffer[1358] = 1358;
 buffer[1359] = 1359;
 buffer[1360] = 1360;
 buffer[1361] = 1361;
 buffer[1362] = 1362;
 buffer[1363] = 1363;
 buffer[1364] = 1364;
 buffer[1365] = 1365;
 buffer[1366] = 1366;
 buffer[1367] = 1367;
 buffer[1368] = 1368;
 buffer[1369] = 1369;
 buffer[1370] = 1370;
 buffer[1371] = 1371;
 buffer[1372] = 1372;
 buffer[1373] = 1373;
 buffer[1374] = 1374;
 buffer[1375] = 1375;
 buffer[1376] = 1376;
 buffer[1377] = 1377;
 buffer[1378] = 1378;
 buffer[1379] = 1379;
 buffer[1380] = 1380;
 buffer[1381] = 1381;
 buffer[1382] = 1382;
 buffer[1383] = 1383;
 buffer[1384] = 1384;
 buffer[1385] = 1385;
 buffer[1386] = 1386;
 buffer[1387] = 1387;
 buffer[1388] = 1388;
 buffer[1389] = 1389;
 buffer[1390] = 1390;
 buffer[1391] = 1391;
 buffer[1392] = 1392;
 buffer[1393] = 1393;
 buffer[1394] = 1394;
 buffer[1395] = 1395;
 buffer[1396] = 1396;
 buffer[1397] = 1397;
 buffer[1398] = 1398;
 buffer[1399] = 1399;
 buffer[1400] = 1400;
 buffer[1401] = 1401;
 buffer[1402] = 1402;
 buffer[1403] = 1403;
 buffer[1404] = 1404;
 buffer[1405] = 1405;
 buffer[1406] = 1406;
 buffer[1407] = 1407;
 buffer[1408] = 1408;
 buffer[1409] = 1409;
 buffer[1410] = 1410;
 buffer[1411] = 1411;
 buffer[1412] = 1412;
 buffer[1413] = 1413;
 buffer[1414] = 1414;
 buffer[1415] = 1415;
 buffer[1416] = 1416;
 buffer[1417] = 1417;
 buffer[1418] = 1418;
 buffer[1419] = 1419;
 buffer[1420] = 1420;
 buffer[1421] = 1421;
 buffer[1422] = 1422;
 buffer[1423] = 1423;
 buffer[1424] = 1424;
 buffer[1425] = 1425;
 buffer[1426] = 1426;
 buffer[1427] = 1427;
 buffer[1428] = 1428;
 buffer[1429] = 1429;
 buffer[1430] = 1430;
 buffer[1431] = 1431;
 buffer[1432] = 1432;
 buffer[1433] = 1433;
 buffer[1434] = 1434;
 buffer[1435] = 1435;
 buffer[1436] = 1436;
 buffer[1437] = 1437;
 buffer[1438] = 1438;
 buffer[1439] = 1439;
 buffer[1440] = 1440;
 buffer[1441] = 1441;
 buffer[1442] = 1442;
 buffer[1443] = 1443;
 buffer[1444] = 1444;
 buffer[1445] = 1445;
 buffer[1446] = 1446;
 buffer[1447] = 1447;
 buffer[1448] = 1448;
 buffer[1449] = 1449;
 buffer[1450] = 1450;
 buffer[1451] = 1451;
 buffer[1452] = 1452;
 buffer[1453] = 1453;
 buffer[1454] = 1454;
 buffer[1455] = 1455;
 buffer[1456] = 1456;
 buffer[1457] = 1457;
 buffer[1458] = 1458;
 buffer[1459] = 1459;
 buffer[1460] = 1460;
 buffer[1461] = 1461;
 buffer[1462] = 1462;
 buffer[1463] = 1463;
 buffer[1464] = 1464;
 buffer[1465] = 1465;
 buffer[1466] = 1466;
 buffer[1467] = 1467;
 buffer[1468] = 1468;
 buffer[1469] = 1469;
 buffer[1470] = 1470;
 buffer[1471] = 1471;
 buffer[1472] = 1472;
 buffer[1473] = 1473;
 buffer[1474] = 1474;
 buffer[1475] = 1475;
 buffer[1476] = 1476;
 buffer[1477] = 1477;
 buffer[1478] = 1478;
 buffer[1479] = 1479;
 buffer[1480] = 1480;
 buffer[1481] = 1481;
 buffer[1482] = 1482;
 buffer[1483] = 1483;
 buffer[1484] = 1484;
 buffer[1485] = 1485;
 buffer[1486] = 1486;
 buffer[1487] = 1487;
 buffer[1488] = 1488;
 buffer[1489] = 1489;
 buffer[1490] = 1490;
 buffer[1491] = 1491;
 buffer[1492] = 1492;
 buffer[1493] = 1493;
 buffer[1494] = 1494;
 buffer[1495] = 1495;
 buffer[1496] = 1496;
 buffer[1497] = 1497;
 buffer[1498] = 1498;
 buffer[1499] = 1499;
 buffer[1500] = 1500;
 buffer[1501] = 1501;
 buffer[1502] = 1502;
 buffer[1503] = 1503;
 buffer[1504] = 1504;
 buffer[1505] = 1505;
 buffer[1506] = 1506;
 buffer[1507] = 1507;
 buffer[1508] = 1508;
 buffer[1509] = 1509;
 buffer[1510] = 1510;
 buffer[1511] = 1511;
 buffer[1512] = 1512;
 buffer[1513] = 1513;
 buffer[1514] = 1514;
 buffer[1515] = 1515;
 buffer[1516] = 1516;
 buffer[1517] = 1517;
 buffer[1518] = 1518;
 buffer[1519] = 1519;
 buffer[1520] = 1520;
 buffer[1521] = 1521;
 buffer[1522] = 1522;
 buffer[1523] = 1523;
 buffer[1524] = 1524;
 buffer[1525] = 1525;
 buffer[1526] = 1526;
 buffer[1527] = 1527;
 buffer[1528] = 1528;
 buffer[1529] = 1529;
 buffer[1530] = 1530;
 buffer[1531] = 1531;
 buffer[1532] = 1532;
 buffer[1533] = 1533;
 buffer[1534] = 1534;
 buffer[1535] = 1535;
 buffer[1536] = 1536;
 buffer[1537] = 1537;
 buffer[1538] = 1538;
 buffer[1539] = 1539;
 buffer[1540] = 1540;
 buffer[1541] = 1541;
 buffer[1542] = 1542;
 buffer[1543] = 1543;
 buffer[1544] = 1544;
 buffer[1545] = 1545;
 buffer[1546] = 1546;
 buffer[1547] = 1547;
 buffer[1548] = 1548;
 buffer[1549] = 1549;
 buffer[1550] = 1550;
 buffer[1551] = 1551;
 buffer[1552] = 1552;
 buffer[1553] = 1553;
 buffer[1554] = 1554;
 buffer[1555] = 1555;
 buffer[1556] = 1556;
 buffer[1557] = 1557;
 buffer[1558] = 1558;
 buffer[1559] = 1559;
 buffer[1560] = 1560;
 buffer[1561] = 1561;
 buffer[1562] = 1562;
 buffer[1563] = 1563;
 buffer[1564] = 1564;
 buffer[1565] = 1565;
 buffer[1566] = 1566;
 buffer[1567] = 1567;
 buffer[1568] = 1568;
 buffer[1569] = 1569;
 buffer[1570] = 1570;
 buffer[1571] = 1571;
 buffer[1572] = 1572;
 buffer[1573] = 1573;
 buffer[1574] = 1574;
 buffer[1575] = 1575;
 buffer[1576] = 1576;
 buffer[1577] = 1577;
 buffer[1578] = 1578;
 buffer[1579] = 1579;
 buffer[1580] = 1580;
 buffer[1581] = 1581;
 buffer[1582] = 1582;
 buffer[1583] = 1583;
 buffer[1584] = 1584;
 buffer[1585] = 1585;
 buffer[1586] = 1586;
 buffer[1587] = 1587;
 buffer[1588] = 1588;
 buffer[1589] = 1589;
 buffer[1590] = 1590;
 buffer[1591] = 1591;
 buffer[1592] = 1592;
 buffer[1593] = 1593;
 buffer[1594] = 1594;
 buffer[1595] = 1595;
 buffer[1596] = 1596;
 buffer[1597] = 1597;
 buffer[1598] = 1598;
 buffer[1599] = 1599;
 buffer[1600] = 1600;
 buffer[1601] = 1601;
 buffer[1602] = 1602;
 buffer[1603] = 1603;
 buffer[1604] = 1604;
 buffer[1605] = 1605;
 buffer[1606] = 1606;
 buffer[1607] = 1607;
 buffer[1608] = 1608;
 buffer[1609] = 1609;
 buffer[1610] = 1610;
 buffer[1611] = 1611;
 buffer[1612] = 1612;
 buffer[1613] = 1613;
 buffer[1614] = 1614;
 buffer[1615] = 1615;
 buffer[1616] = 1616;
 buffer[1617] = 1617;
 buffer[1618] = 1618;
 buffer[1619] = 1619;
 buffer[1620] = 1620;
 buffer[1621] = 1621;
 buffer[1622] = 1622;
 buffer[1623] = 1623;
 buffer[1624] = 1624;
 buffer[1625] = 1625;
 buffer[1626] = 1626;
 buffer[1627] = 1627;
 buffer[1628] = 1628;
 buffer[1629] = 1629;
 buffer[1630] = 1630;
 buffer[1631] = 1631;
 buffer[1632] = 1632;
 buffer[1633] = 1633;
 buffer[1634] = 1634;
 buffer[1635] = 1635;
 buffer[1636] = 1636;
 buffer[1637] = 1637;
 buffer[1638] = 1638;
 buffer[1639] = 1639;
 buffer[1640] = 1640;
 buffer[1641] = 1641;
 buffer[1642] = 1642;
 buffer[1643] = 1643;
 buffer[1644] = 1644;
 buffer[1645] = 1645;
 buffer[1646] = 1646;
 buffer[1647] = 1647;
 buffer[1648] = 1648;
 buffer[1649] = 1649;
 buffer[1650] = 1650;
 buffer[1651] = 1651;
 buffer[1652] = 1652;
 buffer[1653] = 1653;
 buffer[1654] = 1654;
 buffer[1655] = 1655;
 buffer[1656] = 1656;
 buffer[1657] = 1657;
 buffer[1658] = 1658;
 buffer[1659] = 1659;
 buffer[1660] = 1660;
 buffer[1661] = 1661;
 buffer[1662] = 1662;
 buffer[1663] = 1663;
 buffer[1664] = 1664;
 buffer[1665] = 1665;
 buffer[1666] = 1666;
 buffer[1667] = 1667;
 buffer[1668] = 1668;
 buffer[1669] = 1669;
 buffer[1670] = 1670;
 buffer[1671] = 1671;
 buffer[1672] = 1672;
 buffer[1673] = 1673;
 buffer[1674] = 1674;
 buffer[1675] = 1675;
 buffer[1676] = 1676;
 buffer[1677] = 1677;
 buffer[1678] = 1678;
 buffer[1679] = 1679;
 buffer[1680] = 1680;
 buffer[1681] = 1681;
 buffer[1682] = 1682;
 buffer[1683] = 1683;
 buffer[1684] = 1684;
 buffer[1685] = 1685;
 buffer[1686] = 1686;
 buffer[1687] = 1687;
 buffer[1688] = 1688;
 buffer[1689] = 1689;
 buffer[1690] = 1690;
 buffer[1691] = 1691;
 buffer[1692] = 1692;
 buffer[1693] = 1693;
 buffer[1694] = 1694;
 buffer[1695] = 1695;
 buffer[1696] = 1696;
 buffer[1697] = 1697;
 buffer[1698] = 1698;
 buffer[1699] = 1699;
 buffer[1700] = 1700;
 buffer[1701] = 1701;
 buffer[1702] = 1702;
 buffer[1703] = 1703;
 buffer[1704] = 1704;
 buffer[1705] = 1705;
 buffer[1706] = 1706;
 buffer[1707] = 1707;
 buffer[1708] = 1708;
 buffer[1709] = 1709;
 buffer[1710] = 1710;
 buffer[1711] = 1711;
 buffer[1712] = 1712;
 buffer[1713] = 1713;
 buffer[1714] = 1714;
 buffer[1715] = 1715;
 buffer[1716] = 1716;
 buffer[1717] = 1717;
 buffer[1718] = 1718;
 buffer[1719] = 1719;
 buffer[1720] = 1720;
 buffer[1721] = 1721;
 buffer[1722] = 1722;
 buffer[1723] = 1723;
 buffer[1724] = 1724;
 buffer[1725] = 1725;
 buffer[1726] = 1726;
 buffer[1727] = 1727;
 buffer[1728] = 1728;
 buffer[1729] = 1729;
 buffer[1730] = 1730;
 buffer[1731] = 1731;
 buffer[1732] = 1732;
 buffer[1733] = 1733;
 buffer[1734] = 1734;
 buffer[1735] = 1735;
 buffer[1736] = 1736;
 buffer[1737] = 1737;
 buffer[1738] = 1738;
 buffer[1739] = 1739;
 buffer[1740] = 1740;
 buffer[1741] = 1741;
 buffer[1742] = 1742;
 buffer[1743] = 1743;
 buffer[1744] = 1744;
 buffer[1745] = 1745;
 buffer[1746] = 1746;
 buffer[1747] = 1747;
 buffer[1748] = 1748;
 buffer[1749] = 1749;
 buffer[1750] = 1750;
 buffer[1751] = 1751;
 buffer[1752] = 1752;
 buffer[1753] = 1753;
 buffer[1754] = 1754;
 buffer[1755] = 1755;
 buffer[1756] = 1756;
 buffer[1757] = 1757;
 buffer[1758] = 1758;
 buffer[1759] = 1759;
 buffer[1760] = 1760;
 buffer[1761] = 1761;
 buffer[1762] = 1762;
 buffer[1763] = 1763;
 buffer[1764] = 1764;
 buffer[1765] = 1765;
 buffer[1766] = 1766;
 buffer[1767] = 1767;
 buffer[1768] = 1768;
 buffer[1769] = 1769;
 buffer[1770] = 1770;
 buffer[1771] = 1771;
 buffer[1772] = 1772;
 buffer[1773] = 1773;
 buffer[1774] = 1774;
 buffer[1775] = 1775;
 buffer[1776] = 1776;
 buffer[1777] = 1777;
 buffer[1778] = 1778;
 buffer[1779] = 1779;
 buffer[1780] = 1780;
 buffer[1781] = 1781;
 buffer[1782] = 1782;
 buffer[1783] = 1783;
 buffer[1784] = 1784;
 buffer[1785] = 1785;
 buffer[1786] = 1786;
 buffer[1787] = 1787;
 buffer[1788] = 1788;
 buffer[1789] = 1789;
 buffer[1790] = 1790;
 buffer[1791] = 1791;
 buffer[1792] = 1792;
 buffer[1793] = 1793;
 buffer[1794] = 1794;
 buffer[1795] = 1795;
 buffer[1796] = 1796;
 buffer[1797] = 1797;
 buffer[1798] = 1798;
 buffer[1799] = 1799;
 buffer[1800] = 1800;
 buffer[1801] = 1801;
 buffer[1802] = 1802;
 buffer[1803] = 1803;
 buffer[1804] = 1804;
 buffer[1805] = 1805;
 buffer[1806] = 1806;
 buffer[1807] = 1807;
 buffer[1808] = 1808;
 buffer[1809] = 1809;
 buffer[1810] = 1810;
 buffer[1811] = 1811;
 buffer[1812] = 1812;
 buffer[1813] = 1813;
 buffer[1814] = 1814;
 buffer[1815] = 1815;
 buffer[1816] = 1816;
 buffer[1817] = 1817;
 buffer[1818] = 1818;
 buffer[1819] = 1819;
 buffer[1820] = 1820;
 buffer[1821] = 1821;
 buffer[1822] = 1822;
 buffer[1823] = 1823;
 buffer[1824] = 1824;
 buffer[1825] = 1825;
 buffer[1826] = 1826;
 buffer[1827] = 1827;
 buffer[1828] = 1828;
 buffer[1829] = 1829;
 buffer[1830] = 1830;
 buffer[1831] = 1831;
 buffer[1832] = 1832;
 buffer[1833] = 1833;
 buffer[1834] = 1834;
 buffer[1835] = 1835;
 buffer[1836] = 1836;
 buffer[1837] = 1837;
 buffer[1838] = 1838;
 buffer[1839] = 1839;
 buffer[1840] = 1840;
 buffer[1841] = 1841;
 buffer[1842] = 1842;
 buffer[1843] = 1843;
 buffer[1844] = 1844;
 buffer[1845] = 1845;
 buffer[1846] = 1846;
 buffer[1847] = 1847;
 buffer[1848] = 1848;
 buffer[1849] = 1849;
 buffer[1850] = 1850;
 buffer[1851] = 1851;
 buffer[1852] = 1852;
 buffer[1853] = 1853;
 buffer[1854] = 1854;
 buffer[1855] = 1855;
 buffer[1856] = 1856;
 buffer[1857] = 1857;
 buffer[1858] = 1858;
 buffer[1859] = 1859;
 buffer[1860] = 1860;
 buffer[1861] = 1861;
 buffer[1862] = 1862;
 buffer[1863] = 1863;
 buffer[1864] = 1864;
 buffer[1865] = 1865;
 buffer[1866] = 1866;
 buffer[1867] = 1867;
 buffer[1868] = 1868;
 buffer[1869] = 1869;
 buffer[1870] = 1870;
 buffer[1871] = 1871;
 buffer[1872] = 1872;
 buffer[1873] = 1873;
 buffer[1874] = 1874;
 buffer[1875] = 1875;
 buffer[1876] = 1876;
 buffer[1877] = 1877;
 buffer[1878] = 1878;
 buffer[1879] = 1879;
 buffer[1880] = 1880;
 buffer[1881] = 1881;
 buffer[1882] = 1882;
 buffer[1883] = 1883;
 buffer[1884] = 1884;
 buffer[1885] = 1885;
 buffer[1886] = 1886;
 buffer[1887] = 1887;
 buffer[1888] = 1888;
 buffer[1889] = 1889;
 buffer[1890] = 1890;
 buffer[1891] = 1891;
 buffer[1892] = 1892;
 buffer[1893] = 1893;
 buffer[1894] = 1894;
 buffer[1895] = 1895;
 buffer[1896] = 1896;
 buffer[1897] = 1897;
 buffer[1898] = 1898;
 buffer[1899] = 1899;
 buffer[1900] = 1900;
 buffer[1901] = 1901;
 buffer[1902] = 1902;
 buffer[1903] = 1903;
 buffer[1904] = 1904;
 buffer[1905] = 1905;
 buffer[1906] = 1906;
 buffer[1907] = 1907;
 buffer[1908] = 1908;
 buffer[1909] = 1909;
 buffer[1910] = 1910;
 buffer[1911] = 1911;
 buffer[1912] = 1912;
 buffer[1913] = 1913;
 buffer[1914] = 1914;
 buffer[1915] = 1915;
 buffer[1916] = 1916;
 buffer[1917] = 1917;
 buffer[1918] = 1918;
 buffer[1919] = 1919;
 buffer[1920] = 1920;
 buffer[1921] = 1921;
 buffer[1922] = 1922;
 buffer[1923] = 1923;
 buffer[1924] = 1924;
 buffer[1925] = 1925;
 buffer[1926] = 1926;
 buffer[1927] = 1927;
 buffer[1928] = 1928;
 buffer[1929] = 1929;
 buffer[1930] = 1930;
 buffer[1931] = 1931;
 buffer[1932] = 1932;
 buffer[1933] = 1933;
 buffer[1934] = 1934;
 buffer[1935] = 1935;
 buffer[1936] = 1936;
 buffer[1937] = 1937;
 buffer[1938] = 1938;
 buffer[1939] = 1939;
 buffer[1940] = 1940;
 buffer[1941] = 1941;
 buffer[1942] = 1942;
 buffer[1943] = 1943;
 buffer[1944] = 1944;
 buffer[1945] = 1945;
 buffer[1946] = 1946;
 buffer[1947] = 1947;
 buffer[1948] = 1948;
 buffer[1949] = 1949;
 buffer[1950] = 1950;
 buffer[1951] = 1951;
 buffer[1952] = 1952;
 buffer[1953] = 1953;
 buffer[1954] = 1954;
 buffer[1955] = 1955;
 buffer[1956] = 1956;
 buffer[1957] = 1957;
 buffer[1958] = 1958;
 buffer[1959] = 1959;
 buffer[1960] = 1960;
 buffer[1961] = 1961;
 buffer[1962] = 1962;
 buffer[1963] = 1963;
 buffer[1964] = 1964;
 buffer[1965] = 1965;
 buffer[1966] = 1966;
 buffer[1967] = 1967;
 buffer[1968] = 1968;
 buffer[1969] = 1969;
 buffer[1970] = 1970;
 buffer[1971] = 1971;
 buffer[1972] = 1972;
 buffer[1973] = 1973;
 buffer[1974] = 1974;
 buffer[1975] = 1975;
 buffer[1976] = 1976;
 buffer[1977] = 1977;
 buffer[1978] = 1978;
 buffer[1979] = 1979;
 buffer[1980] = 1980;
 buffer[1981] = 1981;
 buffer[1982] = 1982;
 buffer[1983] = 1983;
 buffer[1984] = 1984;
 buffer[1985] = 1985;
 buffer[1986] = 1986;
 buffer[1987] = 1987;
 buffer[1988] = 1988;
 buffer[1989] = 1989;
 buffer[1990] = 1990;
 buffer[1991] = 1991;
 buffer[1992] = 1992;
 buffer[1993] = 1993;
 buffer[1994] = 1994;
 buffer[1995] = 1995;
 buffer[1996] = 1996;
 buffer[1997] = 1997;
 buffer[1998] = 1998;
 buffer[1999] = 1999;
 buffer[2000] = 2000;
 buffer[2001] = 2001;
 buffer[2002] = 2002;
 buffer[2003] = 2003;
 buffer[2004] = 2004;
 buffer[2005] = 2005;
 buffer[2006] = 2006;
 buffer[2007] = 2007;
 buffer[2008] = 2008;
 buffer[2009] = 2009;
 buffer[2010] = 2010;
 buffer[2011] = 2011;
 buffer[2012] = 2012;
 buffer[2013] = 2013;
 buffer[2014] = 2014;
 buffer[2015] = 2015;
 buffer[2016] = 2016;
 buffer[2017] = 2017;
 buffer[2018] = 2018;
 buffer[2019] = 2019;
 buffer[2020] = 2020;
 buffer[2021] = 2021;
 buffer[2022] = 2022;
 buffer[2023] = 2023;
 buffer[2024] = 2024;
 buffer[2025] = 2025;
 buffer[2026] = 2026;
 buffer[2027] = 2027;
 buffer[2028] = 2028;
 buffer[2029] = 2029;
 buffer[2030] = 2030;
 buffer[2031] = 2031;
 buffer[2032] = 2032;
 buffer[2033] = 2033;
 buffer[2034] = 2034;
 buffer[2035] = 2035;
 buffer[2036] = 2036;
 buffer[2037] = 2037;
 buffer[2038] = 2038;
 buffer[2039] = 2039;
 buffer[2040] = 2040;
 buffer[2041] = 2041;
 buffer[2042] = 2042;
 buffer[2043] = 2043;
 buffer[2044] = 2044;
 buffer[2045] = 2045;
 buffer[2046] = 2046;
 buffer[2047] = 2047;
 buffer[2048] = 2048;
 buffer[2049] = 2049;
 buffer[2050] = 2050;
 buffer[2051] = 2051;
 buffer[2052] = 2052;
 buffer[2053] = 2053;
 buffer[2054] = 2054;
 buffer[2055] = 2055;
 buffer[2056] = 2056;
 buffer[2057] = 2057;
 buffer[2058] = 2058;
 buffer[2059] = 2059;
 buffer[2060] = 2060;
 buffer[2061] = 2061;
 buffer[2062] = 2062;
 buffer[2063] = 2063;
 buffer[2064] = 2064;
 buffer[2065] = 2065;
 buffer[2066] = 2066;
 buffer[2067] = 2067;
 buffer[2068] = 2068;
 buffer[2069] = 2069;
 buffer[2070] = 2070;
 buffer[2071] = 2071;
 buffer[2072] = 2072;
 buffer[2073] = 2073;
 buffer[2074] = 2074;
 buffer[2075] = 2075;
 buffer[2076] = 2076;
 buffer[2077] = 2077;
 buffer[2078] = 2078;
 buffer[2079] = 2079;
 buffer[2080] = 2080;
 buffer[2081] = 2081;
 buffer[2082] = 2082;
 buffer[2083] = 2083;
 buffer[2084] = 2084;
 buffer[2085] = 2085;
 buffer[2086] = 2086;
 buffer[2087] = 2087;
 buffer[2088] = 2088;
 buffer[2089] = 2089;
 buffer[2090] = 2090;
 buffer[2091] = 2091;
 buffer[2092] = 2092;
 buffer[2093] = 2093;
 buffer[2094] = 2094;
 buffer[2095] = 2095;
 buffer[2096] = 2096;
 buffer[2097] = 2097;
 buffer[2098] = 2098;
 buffer[2099] = 2099;
 buffer[2100] = 2100;
 buffer[2101] = 2101;
 buffer[2102] = 2102;
 buffer[2103] = 2103;
 buffer[2104] = 2104;
 buffer[2105] = 2105;
 buffer[2106] = 2106;
 buffer[2107] = 2107;
 buffer[2108] = 2108;
 buffer[2109] = 2109;
 buffer[2110] = 2110;
 buffer[2111] = 2111;
 buffer[2112] = 2112;
 buffer[2113] = 2113;
 buffer[2114] = 2114;
 buffer[2115] = 2115;
 buffer[2116] = 2116;
 buffer[2117] = 2117;
 buffer[2118] = 2118;
 buffer[2119] = 2119;
 buffer[2120] = 2120;
 buffer[2121] = 2121;
 buffer[2122] = 2122;
 buffer[2123] = 2123;
 buffer[2124] = 2124;
 buffer[2125] = 2125;
 buffer[2126] = 2126;
 buffer[2127] = 2127;
 buffer[2128] = 2128;
 buffer[2129] = 2129;
 buffer[2130] = 2130;
 buffer[2131] = 2131;
 buffer[2132] = 2132;
 buffer[2133] = 2133;
 buffer[2134] = 2134;
 buffer[2135] = 2135;
 buffer[2136] = 2136;
 buffer[2137] = 2137;
 buffer[2138] = 2138;
 buffer[2139] = 2139;
 buffer[2140] = 2140;
 buffer[2141] = 2141;
 buffer[2142] = 2142;
 buffer[2143] = 2143;
 buffer[2144] = 2144;
 buffer[2145] = 2145;
 buffer[2146] = 2146;
 buffer[2147] = 2147;
 buffer[2148] = 2148;
 buffer[2149] = 2149;
 buffer[2150] = 2150;
 buffer[2151] = 2151;
 buffer[2152] = 2152;
 buffer[2153] = 2153;
 buffer[2154] = 2154;
 buffer[2155] = 2155;
 buffer[2156] = 2156;
 buffer[2157] = 2157;
 buffer[2158] = 2158;
 buffer[2159] = 2159;
 buffer[2160] = 2160;
 buffer[2161] = 2161;
 buffer[2162] = 2162;
 buffer[2163] = 2163;
 buffer[2164] = 2164;
 buffer[2165] = 2165;
 buffer[2166] = 2166;
 buffer[2167] = 2167;
 buffer[2168] = 2168;
 buffer[2169] = 2169;
 buffer[2170] = 2170;
 buffer[2171] = 2171;
 buffer[2172] = 2172;
 buffer[2173] = 2173;
 buffer[2174] = 2174;
 buffer[2175] = 2175;
 buffer[2176] = 2176;
 buffer[2177] = 2177;
 buffer[2178] = 2178;
 buffer[2179] = 2179;
 buffer[2180] = 2180;
 buffer[2181] = 2181;
 buffer[2182] = 2182;
 buffer[2183] = 2183;
 buffer[2184] = 2184;
 buffer[2185] = 2185;
 buffer[2186] = 2186;
 buffer[2187] = 2187;
 buffer[2188] = 2188;
 buffer[2189] = 2189;
 buffer[2190] = 2190;
 buffer[2191] = 2191;
 buffer[2192] = 2192;
 buffer[2193] = 2193;
 buffer[2194] = 2194;
 buffer[2195] = 2195;
 buffer[2196] = 2196;
 buffer[2197] = 2197;
 buffer[2198] = 2198;
 buffer[2199] = 2199;
 buffer[2200] = 2200;
 buffer[2201] = 2201;
 buffer[2202] = 2202;
 buffer[2203] = 2203;
 buffer[2204] = 2204;
 buffer[2205] = 2205;
 buffer[2206] = 2206;
 buffer[2207] = 2207;
 buffer[2208] = 2208;
 buffer[2209] = 2209;
 buffer[2210] = 2210;
 buffer[2211] = 2211;
 buffer[2212] = 2212;
 buffer[2213] = 2213;
 buffer[2214] = 2214;
 buffer[2215] = 2215;
 buffer[2216] = 2216;
 buffer[2217] = 2217;
 buffer[2218] = 2218;
 buffer[2219] = 2219;
 buffer[2220] = 2220;
 buffer[2221] = 2221;
 buffer[2222] = 2222;
 buffer[2223] = 2223;
 buffer[2224] = 2224;
 buffer[2225] = 2225;
 buffer[2226] = 2226;
 buffer[2227] = 2227;
 buffer[2228] = 2228;
 buffer[2229] = 2229;
 buffer[2230] = 2230;
 buffer[2231] = 2231;
 buffer[2232] = 2232;
 buffer[2233] = 2233;
 buffer[2234] = 2234;
 buffer[2235] = 2235;
 buffer[2236] = 2236;
 buffer[2237] = 2237;
 buffer[2238] = 2238;
 buffer[2239] = 2239;
 buffer[2240] = 2240;
 buffer[2241] = 2241;
 buffer[2242] = 2242;
 buffer[2243] = 2243;
 buffer[2244] = 2244;
 buffer[2245] = 2245;
 buffer[2246] = 2246;
 buffer[2247] = 2247;
 buffer[2248] = 2248;
 buffer[2249] = 2249;
 buffer[2250] = 2250;
 buffer[2251] = 2251;
 buffer[2252] = 2252;
 buffer[2253] = 2253;
 buffer[2254] = 2254;
 buffer[2255] = 2255;
 buffer[2256] = 2256;
 buffer[2257] = 2257;
 buffer[2258] = 2258;
 buffer[2259] = 2259;
 buffer[2260] = 2260;
 buffer[2261] = 2261;
 buffer[2262] = 2262;
 buffer[2263] = 2263;
 buffer[2264] = 2264;
 buffer[2265] = 2265;
 buffer[2266] = 2266;
 buffer[2267] = 2267;
 buffer[2268] = 2268;
 buffer[2269] = 2269;
 buffer[2270] = 2270;
 buffer[2271] = 2271;
 buffer[2272] = 2272;
 buffer[2273] = 2273;
 buffer[2274] = 2274;
 buffer[2275] = 2275;
 buffer[2276] = 2276;
 buffer[2277] = 2277;
 buffer[2278] = 2278;
 buffer[2279] = 2279;
 buffer[2280] = 2280;
 buffer[2281] = 2281;
 buffer[2282] = 2282;
 buffer[2283] = 2283;
 buffer[2284] = 2284;
 buffer[2285] = 2285;
 buffer[2286] = 2286;
 buffer[2287] = 2287;
 buffer[2288] = 2288;
 buffer[2289] = 2289;
 buffer[2290] = 2290;
 buffer[2291] = 2291;
 buffer[2292] = 2292;
 buffer[2293] = 2293;
 buffer[2294] = 2294;
 buffer[2295] = 2295;
 buffer[2296] = 2296;
 buffer[2297] = 2297;
 buffer[2298] = 2298;
 buffer[2299] = 2299;
 buffer[2300] = 2300;
 buffer[2301] = 2301;
 buffer[2302] = 2302;
 buffer[2303] = 2303;
 buffer[2304] = 2304;
 buffer[2305] = 2305;
 buffer[2306] = 2306;
 buffer[2307] = 2307;
 buffer[2308] = 2308;
 buffer[2309] = 2309;
 buffer[2310] = 2310;
 buffer[2311] = 2311;
 buffer[2312] = 2312;
 buffer[2313] = 2313;
 buffer[2314] = 2314;
 buffer[2315] = 2315;
 buffer[2316] = 2316;
 buffer[2317] = 2317;
 buffer[2318] = 2318;
 buffer[2319] = 2319;
 buffer[2320] = 2320;
 buffer[2321] = 2321;
 buffer[2322] = 2322;
 buffer[2323] = 2323;
 buffer[2324] = 2324;
 buffer[2325] = 2325;
 buffer[2326] = 2326;
 buffer[2327] = 2327;
 buffer[2328] = 2328;
 buffer[2329] = 2329;
 buffer[2330] = 2330;
 buffer[2331] = 2331;
 buffer[2332] = 2332;
 buffer[2333] = 2333;
 buffer[2334] = 2334;
 buffer[2335] = 2335;
 buffer[2336] = 2336;
 buffer[2337] = 2337;
 buffer[2338] = 2338;
 buffer[2339] = 2339;
 buffer[2340] = 2340;
 buffer[2341] = 2341;
 buffer[2342] = 2342;
 buffer[2343] = 2343;
 buffer[2344] = 2344;
 buffer[2345] = 2345;
 buffer[2346] = 2346;
 buffer[2347] = 2347;
 buffer[2348] = 2348;
 buffer[2349] = 2349;
 buffer[2350] = 2350;
 buffer[2351] = 2351;
 buffer[2352] = 2352;
 buffer[2353] = 2353;
 buffer[2354] = 2354;
 buffer[2355] = 2355;
 buffer[2356] = 2356;
 buffer[2357] = 2357;
 buffer[2358] = 2358;
 buffer[2359] = 2359;
 buffer[2360] = 2360;
 buffer[2361] = 2361;
 buffer[2362] = 2362;
 buffer[2363] = 2363;
 buffer[2364] = 2364;
 buffer[2365] = 2365;
 buffer[2366] = 2366;
 buffer[2367] = 2367;
 buffer[2368] = 2368;
 buffer[2369] = 2369;
 buffer[2370] = 2370;
 buffer[2371] = 2371;
 buffer[2372] = 2372;
 buffer[2373] = 2373;
 buffer[2374] = 2374;
 buffer[2375] = 2375;
 buffer[2376] = 2376;
 buffer[2377] = 2377;
 buffer[2378] = 2378;
 buffer[2379] = 2379;
 buffer[2380] = 2380;
 buffer[2381] = 2381;
 buffer[2382] = 2382;
 buffer[2383] = 2383;
 buffer[2384] = 2384;
 buffer[2385] = 2385;
 buffer[2386] = 2386;
 buffer[2387] = 2387;
 buffer[2388] = 2388;
 buffer[2389] = 2389;
 buffer[2390] = 2390;
 buffer[2391] = 2391;
 buffer[2392] = 2392;
 buffer[2393] = 2393;
 buffer[2394] = 2394;
 buffer[2395] = 2395;
 buffer[2396] = 2396;
 buffer[2397] = 2397;
 buffer[2398] = 2398;
 buffer[2399] = 2399;
end

endmodule

module M_multiplex_display_mem_background(
input      [0:0]             in_background_wenable0,
input       [7:0]     in_background_wdata0,
input      [11:0]                in_background_addr0,
input      [0:0]             in_background_wenable1,
input      [7:0]                 in_background_wdata1,
input      [11:0]                in_background_addr1,
output reg  [7:0]     out_background_rdata0,
output reg  [7:0]     out_background_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2399:0];
always @(posedge clock0) begin
  if (in_background_wenable0) begin
    buffer[in_background_addr0] <= in_background_wdata0;
  end else begin
    out_background_rdata0 <= buffer[in_background_addr0];
  end
end
always @(posedge clock1) begin
  if (in_background_wenable1) begin
    buffer[in_background_addr1] <= in_background_wdata1;
  end else begin
    out_background_rdata1 <= buffer[in_background_addr1];
  end
end
initial begin
 buffer[0] = 2399;
 buffer[1] = 2398;
 buffer[2] = 2397;
 buffer[3] = 2396;
 buffer[4] = 2395;
 buffer[5] = 2394;
 buffer[6] = 2393;
 buffer[7] = 2392;
 buffer[8] = 2391;
 buffer[9] = 2390;
 buffer[10] = 2389;
 buffer[11] = 2388;
 buffer[12] = 2387;
 buffer[13] = 2386;
 buffer[14] = 2385;
 buffer[15] = 2384;
 buffer[16] = 2383;
 buffer[17] = 2382;
 buffer[18] = 2381;
 buffer[19] = 2380;
 buffer[20] = 2379;
 buffer[21] = 2378;
 buffer[22] = 2377;
 buffer[23] = 2376;
 buffer[24] = 2375;
 buffer[25] = 2374;
 buffer[26] = 2373;
 buffer[27] = 2372;
 buffer[28] = 2371;
 buffer[29] = 2370;
 buffer[30] = 2369;
 buffer[31] = 2368;
 buffer[32] = 2367;
 buffer[33] = 2366;
 buffer[34] = 2365;
 buffer[35] = 2364;
 buffer[36] = 2363;
 buffer[37] = 2362;
 buffer[38] = 2361;
 buffer[39] = 2360;
 buffer[40] = 2359;
 buffer[41] = 2358;
 buffer[42] = 2357;
 buffer[43] = 2356;
 buffer[44] = 2355;
 buffer[45] = 2354;
 buffer[46] = 2353;
 buffer[47] = 2352;
 buffer[48] = 2351;
 buffer[49] = 2350;
 buffer[50] = 2349;
 buffer[51] = 2348;
 buffer[52] = 2347;
 buffer[53] = 2346;
 buffer[54] = 2345;
 buffer[55] = 2344;
 buffer[56] = 2343;
 buffer[57] = 2342;
 buffer[58] = 2341;
 buffer[59] = 2340;
 buffer[60] = 2339;
 buffer[61] = 2338;
 buffer[62] = 2337;
 buffer[63] = 2336;
 buffer[64] = 2335;
 buffer[65] = 2334;
 buffer[66] = 2333;
 buffer[67] = 2332;
 buffer[68] = 2331;
 buffer[69] = 2330;
 buffer[70] = 2329;
 buffer[71] = 2328;
 buffer[72] = 2327;
 buffer[73] = 2326;
 buffer[74] = 2325;
 buffer[75] = 2324;
 buffer[76] = 2323;
 buffer[77] = 2322;
 buffer[78] = 2321;
 buffer[79] = 2320;
 buffer[80] = 2319;
 buffer[81] = 2318;
 buffer[82] = 2317;
 buffer[83] = 2316;
 buffer[84] = 2315;
 buffer[85] = 2314;
 buffer[86] = 2313;
 buffer[87] = 2312;
 buffer[88] = 2311;
 buffer[89] = 2310;
 buffer[90] = 2309;
 buffer[91] = 2308;
 buffer[92] = 2307;
 buffer[93] = 2306;
 buffer[94] = 2305;
 buffer[95] = 2304;
 buffer[96] = 2303;
 buffer[97] = 2302;
 buffer[98] = 2301;
 buffer[99] = 2300;
 buffer[100] = 2299;
 buffer[101] = 2298;
 buffer[102] = 2297;
 buffer[103] = 2296;
 buffer[104] = 2295;
 buffer[105] = 2294;
 buffer[106] = 2293;
 buffer[107] = 2292;
 buffer[108] = 2291;
 buffer[109] = 2290;
 buffer[110] = 2289;
 buffer[111] = 2288;
 buffer[112] = 2287;
 buffer[113] = 2286;
 buffer[114] = 2285;
 buffer[115] = 2284;
 buffer[116] = 2283;
 buffer[117] = 2282;
 buffer[118] = 2281;
 buffer[119] = 2280;
 buffer[120] = 2279;
 buffer[121] = 2278;
 buffer[122] = 2277;
 buffer[123] = 2276;
 buffer[124] = 2275;
 buffer[125] = 2274;
 buffer[126] = 2273;
 buffer[127] = 2272;
 buffer[128] = 2271;
 buffer[129] = 2270;
 buffer[130] = 2269;
 buffer[131] = 2268;
 buffer[132] = 2267;
 buffer[133] = 2266;
 buffer[134] = 2265;
 buffer[135] = 2264;
 buffer[136] = 2263;
 buffer[137] = 2262;
 buffer[138] = 2261;
 buffer[139] = 2260;
 buffer[140] = 2259;
 buffer[141] = 2258;
 buffer[142] = 2257;
 buffer[143] = 2256;
 buffer[144] = 2255;
 buffer[145] = 2254;
 buffer[146] = 2253;
 buffer[147] = 2252;
 buffer[148] = 2251;
 buffer[149] = 2250;
 buffer[150] = 2249;
 buffer[151] = 2248;
 buffer[152] = 2247;
 buffer[153] = 2246;
 buffer[154] = 2245;
 buffer[155] = 2244;
 buffer[156] = 2243;
 buffer[157] = 2242;
 buffer[158] = 2241;
 buffer[159] = 2240;
 buffer[160] = 2239;
 buffer[161] = 2238;
 buffer[162] = 2237;
 buffer[163] = 2236;
 buffer[164] = 2235;
 buffer[165] = 2234;
 buffer[166] = 2233;
 buffer[167] = 2232;
 buffer[168] = 2231;
 buffer[169] = 2230;
 buffer[170] = 2229;
 buffer[171] = 2228;
 buffer[172] = 2227;
 buffer[173] = 2226;
 buffer[174] = 2225;
 buffer[175] = 2224;
 buffer[176] = 2223;
 buffer[177] = 2222;
 buffer[178] = 2221;
 buffer[179] = 2220;
 buffer[180] = 2219;
 buffer[181] = 2218;
 buffer[182] = 2217;
 buffer[183] = 2216;
 buffer[184] = 2215;
 buffer[185] = 2214;
 buffer[186] = 2213;
 buffer[187] = 2212;
 buffer[188] = 2211;
 buffer[189] = 2210;
 buffer[190] = 2209;
 buffer[191] = 2208;
 buffer[192] = 2207;
 buffer[193] = 2206;
 buffer[194] = 2205;
 buffer[195] = 2204;
 buffer[196] = 2203;
 buffer[197] = 2202;
 buffer[198] = 2201;
 buffer[199] = 2200;
 buffer[200] = 2199;
 buffer[201] = 2198;
 buffer[202] = 2197;
 buffer[203] = 2196;
 buffer[204] = 2195;
 buffer[205] = 2194;
 buffer[206] = 2193;
 buffer[207] = 2192;
 buffer[208] = 2191;
 buffer[209] = 2190;
 buffer[210] = 2189;
 buffer[211] = 2188;
 buffer[212] = 2187;
 buffer[213] = 2186;
 buffer[214] = 2185;
 buffer[215] = 2184;
 buffer[216] = 2183;
 buffer[217] = 2182;
 buffer[218] = 2181;
 buffer[219] = 2180;
 buffer[220] = 2179;
 buffer[221] = 2178;
 buffer[222] = 2177;
 buffer[223] = 2176;
 buffer[224] = 2175;
 buffer[225] = 2174;
 buffer[226] = 2173;
 buffer[227] = 2172;
 buffer[228] = 2171;
 buffer[229] = 2170;
 buffer[230] = 2169;
 buffer[231] = 2168;
 buffer[232] = 2167;
 buffer[233] = 2166;
 buffer[234] = 2165;
 buffer[235] = 2164;
 buffer[236] = 2163;
 buffer[237] = 2162;
 buffer[238] = 2161;
 buffer[239] = 2160;
 buffer[240] = 2159;
 buffer[241] = 2158;
 buffer[242] = 2157;
 buffer[243] = 2156;
 buffer[244] = 2155;
 buffer[245] = 2154;
 buffer[246] = 2153;
 buffer[247] = 2152;
 buffer[248] = 2151;
 buffer[249] = 2150;
 buffer[250] = 2149;
 buffer[251] = 2148;
 buffer[252] = 2147;
 buffer[253] = 2146;
 buffer[254] = 2145;
 buffer[255] = 2144;
 buffer[256] = 2143;
 buffer[257] = 2142;
 buffer[258] = 2141;
 buffer[259] = 2140;
 buffer[260] = 2139;
 buffer[261] = 2138;
 buffer[262] = 2137;
 buffer[263] = 2136;
 buffer[264] = 2135;
 buffer[265] = 2134;
 buffer[266] = 2133;
 buffer[267] = 2132;
 buffer[268] = 2131;
 buffer[269] = 2130;
 buffer[270] = 2129;
 buffer[271] = 2128;
 buffer[272] = 2127;
 buffer[273] = 2126;
 buffer[274] = 2125;
 buffer[275] = 2124;
 buffer[276] = 2123;
 buffer[277] = 2122;
 buffer[278] = 2121;
 buffer[279] = 2120;
 buffer[280] = 2119;
 buffer[281] = 2118;
 buffer[282] = 2117;
 buffer[283] = 2116;
 buffer[284] = 2115;
 buffer[285] = 2114;
 buffer[286] = 2113;
 buffer[287] = 2112;
 buffer[288] = 2111;
 buffer[289] = 2110;
 buffer[290] = 2109;
 buffer[291] = 2108;
 buffer[292] = 2107;
 buffer[293] = 2106;
 buffer[294] = 2105;
 buffer[295] = 2104;
 buffer[296] = 2103;
 buffer[297] = 2102;
 buffer[298] = 2101;
 buffer[299] = 2100;
 buffer[300] = 2099;
 buffer[301] = 2098;
 buffer[302] = 2097;
 buffer[303] = 2096;
 buffer[304] = 2095;
 buffer[305] = 2094;
 buffer[306] = 2093;
 buffer[307] = 2092;
 buffer[308] = 2091;
 buffer[309] = 2090;
 buffer[310] = 2089;
 buffer[311] = 2088;
 buffer[312] = 2087;
 buffer[313] = 2086;
 buffer[314] = 2085;
 buffer[315] = 2084;
 buffer[316] = 2083;
 buffer[317] = 2082;
 buffer[318] = 2081;
 buffer[319] = 2080;
 buffer[320] = 2079;
 buffer[321] = 2078;
 buffer[322] = 2077;
 buffer[323] = 2076;
 buffer[324] = 2075;
 buffer[325] = 2074;
 buffer[326] = 2073;
 buffer[327] = 2072;
 buffer[328] = 2071;
 buffer[329] = 2070;
 buffer[330] = 2069;
 buffer[331] = 2068;
 buffer[332] = 2067;
 buffer[333] = 2066;
 buffer[334] = 2065;
 buffer[335] = 2064;
 buffer[336] = 2063;
 buffer[337] = 2062;
 buffer[338] = 2061;
 buffer[339] = 2060;
 buffer[340] = 2059;
 buffer[341] = 2058;
 buffer[342] = 2057;
 buffer[343] = 2056;
 buffer[344] = 2055;
 buffer[345] = 2054;
 buffer[346] = 2053;
 buffer[347] = 2052;
 buffer[348] = 2051;
 buffer[349] = 2050;
 buffer[350] = 2049;
 buffer[351] = 2048;
 buffer[352] = 2047;
 buffer[353] = 2046;
 buffer[354] = 2045;
 buffer[355] = 2044;
 buffer[356] = 2043;
 buffer[357] = 2042;
 buffer[358] = 2041;
 buffer[359] = 2040;
 buffer[360] = 2039;
 buffer[361] = 2038;
 buffer[362] = 2037;
 buffer[363] = 2036;
 buffer[364] = 2035;
 buffer[365] = 2034;
 buffer[366] = 2033;
 buffer[367] = 2032;
 buffer[368] = 2031;
 buffer[369] = 2030;
 buffer[370] = 2029;
 buffer[371] = 2028;
 buffer[372] = 2027;
 buffer[373] = 2026;
 buffer[374] = 2025;
 buffer[375] = 2024;
 buffer[376] = 2023;
 buffer[377] = 2022;
 buffer[378] = 2021;
 buffer[379] = 2020;
 buffer[380] = 2019;
 buffer[381] = 2018;
 buffer[382] = 2017;
 buffer[383] = 2016;
 buffer[384] = 2015;
 buffer[385] = 2014;
 buffer[386] = 2013;
 buffer[387] = 2012;
 buffer[388] = 2011;
 buffer[389] = 2010;
 buffer[390] = 2009;
 buffer[391] = 2008;
 buffer[392] = 2007;
 buffer[393] = 2006;
 buffer[394] = 2005;
 buffer[395] = 2004;
 buffer[396] = 2003;
 buffer[397] = 2002;
 buffer[398] = 2001;
 buffer[399] = 2000;
 buffer[400] = 1999;
 buffer[401] = 1998;
 buffer[402] = 1997;
 buffer[403] = 1996;
 buffer[404] = 1995;
 buffer[405] = 1994;
 buffer[406] = 1993;
 buffer[407] = 1992;
 buffer[408] = 1991;
 buffer[409] = 1990;
 buffer[410] = 1989;
 buffer[411] = 1988;
 buffer[412] = 1987;
 buffer[413] = 1986;
 buffer[414] = 1985;
 buffer[415] = 1984;
 buffer[416] = 1983;
 buffer[417] = 1982;
 buffer[418] = 1981;
 buffer[419] = 1980;
 buffer[420] = 1979;
 buffer[421] = 1978;
 buffer[422] = 1977;
 buffer[423] = 1976;
 buffer[424] = 1975;
 buffer[425] = 1974;
 buffer[426] = 1973;
 buffer[427] = 1972;
 buffer[428] = 1971;
 buffer[429] = 1970;
 buffer[430] = 1969;
 buffer[431] = 1968;
 buffer[432] = 1967;
 buffer[433] = 1966;
 buffer[434] = 1965;
 buffer[435] = 1964;
 buffer[436] = 1963;
 buffer[437] = 1962;
 buffer[438] = 1961;
 buffer[439] = 1960;
 buffer[440] = 1959;
 buffer[441] = 1958;
 buffer[442] = 1957;
 buffer[443] = 1956;
 buffer[444] = 1955;
 buffer[445] = 1954;
 buffer[446] = 1953;
 buffer[447] = 1952;
 buffer[448] = 1951;
 buffer[449] = 1950;
 buffer[450] = 1949;
 buffer[451] = 1948;
 buffer[452] = 1947;
 buffer[453] = 1946;
 buffer[454] = 1945;
 buffer[455] = 1944;
 buffer[456] = 1943;
 buffer[457] = 1942;
 buffer[458] = 1941;
 buffer[459] = 1940;
 buffer[460] = 1939;
 buffer[461] = 1938;
 buffer[462] = 1937;
 buffer[463] = 1936;
 buffer[464] = 1935;
 buffer[465] = 1934;
 buffer[466] = 1933;
 buffer[467] = 1932;
 buffer[468] = 1931;
 buffer[469] = 1930;
 buffer[470] = 1929;
 buffer[471] = 1928;
 buffer[472] = 1927;
 buffer[473] = 1926;
 buffer[474] = 1925;
 buffer[475] = 1924;
 buffer[476] = 1923;
 buffer[477] = 1922;
 buffer[478] = 1921;
 buffer[479] = 1920;
 buffer[480] = 1919;
 buffer[481] = 1918;
 buffer[482] = 1917;
 buffer[483] = 1916;
 buffer[484] = 1915;
 buffer[485] = 1914;
 buffer[486] = 1913;
 buffer[487] = 1912;
 buffer[488] = 1911;
 buffer[489] = 1910;
 buffer[490] = 1909;
 buffer[491] = 1908;
 buffer[492] = 1907;
 buffer[493] = 1906;
 buffer[494] = 1905;
 buffer[495] = 1904;
 buffer[496] = 1903;
 buffer[497] = 1902;
 buffer[498] = 1901;
 buffer[499] = 1900;
 buffer[500] = 1899;
 buffer[501] = 1898;
 buffer[502] = 1897;
 buffer[503] = 1896;
 buffer[504] = 1895;
 buffer[505] = 1894;
 buffer[506] = 1893;
 buffer[507] = 1892;
 buffer[508] = 1891;
 buffer[509] = 1890;
 buffer[510] = 1889;
 buffer[511] = 1888;
 buffer[512] = 1887;
 buffer[513] = 1886;
 buffer[514] = 1885;
 buffer[515] = 1884;
 buffer[516] = 1883;
 buffer[517] = 1882;
 buffer[518] = 1881;
 buffer[519] = 1880;
 buffer[520] = 1879;
 buffer[521] = 1878;
 buffer[522] = 1877;
 buffer[523] = 1876;
 buffer[524] = 1875;
 buffer[525] = 1874;
 buffer[526] = 1873;
 buffer[527] = 1872;
 buffer[528] = 1871;
 buffer[529] = 1870;
 buffer[530] = 1869;
 buffer[531] = 1868;
 buffer[532] = 1867;
 buffer[533] = 1866;
 buffer[534] = 1865;
 buffer[535] = 1864;
 buffer[536] = 1863;
 buffer[537] = 1862;
 buffer[538] = 1861;
 buffer[539] = 1860;
 buffer[540] = 1859;
 buffer[541] = 1858;
 buffer[542] = 1857;
 buffer[543] = 1856;
 buffer[544] = 1855;
 buffer[545] = 1854;
 buffer[546] = 1853;
 buffer[547] = 1852;
 buffer[548] = 1851;
 buffer[549] = 1850;
 buffer[550] = 1849;
 buffer[551] = 1848;
 buffer[552] = 1847;
 buffer[553] = 1846;
 buffer[554] = 1845;
 buffer[555] = 1844;
 buffer[556] = 1843;
 buffer[557] = 1842;
 buffer[558] = 1841;
 buffer[559] = 1840;
 buffer[560] = 1839;
 buffer[561] = 1838;
 buffer[562] = 1837;
 buffer[563] = 1836;
 buffer[564] = 1835;
 buffer[565] = 1834;
 buffer[566] = 1833;
 buffer[567] = 1832;
 buffer[568] = 1831;
 buffer[569] = 1830;
 buffer[570] = 1829;
 buffer[571] = 1828;
 buffer[572] = 1827;
 buffer[573] = 1826;
 buffer[574] = 1825;
 buffer[575] = 1824;
 buffer[576] = 1823;
 buffer[577] = 1822;
 buffer[578] = 1821;
 buffer[579] = 1820;
 buffer[580] = 1819;
 buffer[581] = 1818;
 buffer[582] = 1817;
 buffer[583] = 1816;
 buffer[584] = 1815;
 buffer[585] = 1814;
 buffer[586] = 1813;
 buffer[587] = 1812;
 buffer[588] = 1811;
 buffer[589] = 1810;
 buffer[590] = 1809;
 buffer[591] = 1808;
 buffer[592] = 1807;
 buffer[593] = 1806;
 buffer[594] = 1805;
 buffer[595] = 1804;
 buffer[596] = 1803;
 buffer[597] = 1802;
 buffer[598] = 1801;
 buffer[599] = 1800;
 buffer[600] = 1799;
 buffer[601] = 1798;
 buffer[602] = 1797;
 buffer[603] = 1796;
 buffer[604] = 1795;
 buffer[605] = 1794;
 buffer[606] = 1793;
 buffer[607] = 1792;
 buffer[608] = 1791;
 buffer[609] = 1790;
 buffer[610] = 1789;
 buffer[611] = 1788;
 buffer[612] = 1787;
 buffer[613] = 1786;
 buffer[614] = 1785;
 buffer[615] = 1784;
 buffer[616] = 1783;
 buffer[617] = 1782;
 buffer[618] = 1781;
 buffer[619] = 1780;
 buffer[620] = 1779;
 buffer[621] = 1778;
 buffer[622] = 1777;
 buffer[623] = 1776;
 buffer[624] = 1775;
 buffer[625] = 1774;
 buffer[626] = 1773;
 buffer[627] = 1772;
 buffer[628] = 1771;
 buffer[629] = 1770;
 buffer[630] = 1769;
 buffer[631] = 1768;
 buffer[632] = 1767;
 buffer[633] = 1766;
 buffer[634] = 1765;
 buffer[635] = 1764;
 buffer[636] = 1763;
 buffer[637] = 1762;
 buffer[638] = 1761;
 buffer[639] = 1760;
 buffer[640] = 1759;
 buffer[641] = 1758;
 buffer[642] = 1757;
 buffer[643] = 1756;
 buffer[644] = 1755;
 buffer[645] = 1754;
 buffer[646] = 1753;
 buffer[647] = 1752;
 buffer[648] = 1751;
 buffer[649] = 1750;
 buffer[650] = 1749;
 buffer[651] = 1748;
 buffer[652] = 1747;
 buffer[653] = 1746;
 buffer[654] = 1745;
 buffer[655] = 1744;
 buffer[656] = 1743;
 buffer[657] = 1742;
 buffer[658] = 1741;
 buffer[659] = 1740;
 buffer[660] = 1739;
 buffer[661] = 1738;
 buffer[662] = 1737;
 buffer[663] = 1736;
 buffer[664] = 1735;
 buffer[665] = 1734;
 buffer[666] = 1733;
 buffer[667] = 1732;
 buffer[668] = 1731;
 buffer[669] = 1730;
 buffer[670] = 1729;
 buffer[671] = 1728;
 buffer[672] = 1727;
 buffer[673] = 1726;
 buffer[674] = 1725;
 buffer[675] = 1724;
 buffer[676] = 1723;
 buffer[677] = 1722;
 buffer[678] = 1721;
 buffer[679] = 1720;
 buffer[680] = 1719;
 buffer[681] = 1718;
 buffer[682] = 1717;
 buffer[683] = 1716;
 buffer[684] = 1715;
 buffer[685] = 1714;
 buffer[686] = 1713;
 buffer[687] = 1712;
 buffer[688] = 1711;
 buffer[689] = 1710;
 buffer[690] = 1709;
 buffer[691] = 1708;
 buffer[692] = 1707;
 buffer[693] = 1706;
 buffer[694] = 1705;
 buffer[695] = 1704;
 buffer[696] = 1703;
 buffer[697] = 1702;
 buffer[698] = 1701;
 buffer[699] = 1700;
 buffer[700] = 1699;
 buffer[701] = 1698;
 buffer[702] = 1697;
 buffer[703] = 1696;
 buffer[704] = 1695;
 buffer[705] = 1694;
 buffer[706] = 1693;
 buffer[707] = 1692;
 buffer[708] = 1691;
 buffer[709] = 1690;
 buffer[710] = 1689;
 buffer[711] = 1688;
 buffer[712] = 1687;
 buffer[713] = 1686;
 buffer[714] = 1685;
 buffer[715] = 1684;
 buffer[716] = 1683;
 buffer[717] = 1682;
 buffer[718] = 1681;
 buffer[719] = 1680;
 buffer[720] = 1679;
 buffer[721] = 1678;
 buffer[722] = 1677;
 buffer[723] = 1676;
 buffer[724] = 1675;
 buffer[725] = 1674;
 buffer[726] = 1673;
 buffer[727] = 1672;
 buffer[728] = 1671;
 buffer[729] = 1670;
 buffer[730] = 1669;
 buffer[731] = 1668;
 buffer[732] = 1667;
 buffer[733] = 1666;
 buffer[734] = 1665;
 buffer[735] = 1664;
 buffer[736] = 1663;
 buffer[737] = 1662;
 buffer[738] = 1661;
 buffer[739] = 1660;
 buffer[740] = 1659;
 buffer[741] = 1658;
 buffer[742] = 1657;
 buffer[743] = 1656;
 buffer[744] = 1655;
 buffer[745] = 1654;
 buffer[746] = 1653;
 buffer[747] = 1652;
 buffer[748] = 1651;
 buffer[749] = 1650;
 buffer[750] = 1649;
 buffer[751] = 1648;
 buffer[752] = 1647;
 buffer[753] = 1646;
 buffer[754] = 1645;
 buffer[755] = 1644;
 buffer[756] = 1643;
 buffer[757] = 1642;
 buffer[758] = 1641;
 buffer[759] = 1640;
 buffer[760] = 1639;
 buffer[761] = 1638;
 buffer[762] = 1637;
 buffer[763] = 1636;
 buffer[764] = 1635;
 buffer[765] = 1634;
 buffer[766] = 1633;
 buffer[767] = 1632;
 buffer[768] = 1631;
 buffer[769] = 1630;
 buffer[770] = 1629;
 buffer[771] = 1628;
 buffer[772] = 1627;
 buffer[773] = 1626;
 buffer[774] = 1625;
 buffer[775] = 1624;
 buffer[776] = 1623;
 buffer[777] = 1622;
 buffer[778] = 1621;
 buffer[779] = 1620;
 buffer[780] = 1619;
 buffer[781] = 1618;
 buffer[782] = 1617;
 buffer[783] = 1616;
 buffer[784] = 1615;
 buffer[785] = 1614;
 buffer[786] = 1613;
 buffer[787] = 1612;
 buffer[788] = 1611;
 buffer[789] = 1610;
 buffer[790] = 1609;
 buffer[791] = 1608;
 buffer[792] = 1607;
 buffer[793] = 1606;
 buffer[794] = 1605;
 buffer[795] = 1604;
 buffer[796] = 1603;
 buffer[797] = 1602;
 buffer[798] = 1601;
 buffer[799] = 1600;
 buffer[800] = 1599;
 buffer[801] = 1598;
 buffer[802] = 1597;
 buffer[803] = 1596;
 buffer[804] = 1595;
 buffer[805] = 1594;
 buffer[806] = 1593;
 buffer[807] = 1592;
 buffer[808] = 1591;
 buffer[809] = 1590;
 buffer[810] = 1589;
 buffer[811] = 1588;
 buffer[812] = 1587;
 buffer[813] = 1586;
 buffer[814] = 1585;
 buffer[815] = 1584;
 buffer[816] = 1583;
 buffer[817] = 1582;
 buffer[818] = 1581;
 buffer[819] = 1580;
 buffer[820] = 1579;
 buffer[821] = 1578;
 buffer[822] = 1577;
 buffer[823] = 1576;
 buffer[824] = 1575;
 buffer[825] = 1574;
 buffer[826] = 1573;
 buffer[827] = 1572;
 buffer[828] = 1571;
 buffer[829] = 1570;
 buffer[830] = 1569;
 buffer[831] = 1568;
 buffer[832] = 1567;
 buffer[833] = 1566;
 buffer[834] = 1565;
 buffer[835] = 1564;
 buffer[836] = 1563;
 buffer[837] = 1562;
 buffer[838] = 1561;
 buffer[839] = 1560;
 buffer[840] = 1559;
 buffer[841] = 1558;
 buffer[842] = 1557;
 buffer[843] = 1556;
 buffer[844] = 1555;
 buffer[845] = 1554;
 buffer[846] = 1553;
 buffer[847] = 1552;
 buffer[848] = 1551;
 buffer[849] = 1550;
 buffer[850] = 1549;
 buffer[851] = 1548;
 buffer[852] = 1547;
 buffer[853] = 1546;
 buffer[854] = 1545;
 buffer[855] = 1544;
 buffer[856] = 1543;
 buffer[857] = 1542;
 buffer[858] = 1541;
 buffer[859] = 1540;
 buffer[860] = 1539;
 buffer[861] = 1538;
 buffer[862] = 1537;
 buffer[863] = 1536;
 buffer[864] = 1535;
 buffer[865] = 1534;
 buffer[866] = 1533;
 buffer[867] = 1532;
 buffer[868] = 1531;
 buffer[869] = 1530;
 buffer[870] = 1529;
 buffer[871] = 1528;
 buffer[872] = 1527;
 buffer[873] = 1526;
 buffer[874] = 1525;
 buffer[875] = 1524;
 buffer[876] = 1523;
 buffer[877] = 1522;
 buffer[878] = 1521;
 buffer[879] = 1520;
 buffer[880] = 1519;
 buffer[881] = 1518;
 buffer[882] = 1517;
 buffer[883] = 1516;
 buffer[884] = 1515;
 buffer[885] = 1514;
 buffer[886] = 1513;
 buffer[887] = 1512;
 buffer[888] = 1511;
 buffer[889] = 1510;
 buffer[890] = 1509;
 buffer[891] = 1508;
 buffer[892] = 1507;
 buffer[893] = 1506;
 buffer[894] = 1505;
 buffer[895] = 1504;
 buffer[896] = 1503;
 buffer[897] = 1502;
 buffer[898] = 1501;
 buffer[899] = 1500;
 buffer[900] = 1499;
 buffer[901] = 1498;
 buffer[902] = 1497;
 buffer[903] = 1496;
 buffer[904] = 1495;
 buffer[905] = 1494;
 buffer[906] = 1493;
 buffer[907] = 1492;
 buffer[908] = 1491;
 buffer[909] = 1490;
 buffer[910] = 1489;
 buffer[911] = 1488;
 buffer[912] = 1487;
 buffer[913] = 1486;
 buffer[914] = 1485;
 buffer[915] = 1484;
 buffer[916] = 1483;
 buffer[917] = 1482;
 buffer[918] = 1481;
 buffer[919] = 1480;
 buffer[920] = 1479;
 buffer[921] = 1478;
 buffer[922] = 1477;
 buffer[923] = 1476;
 buffer[924] = 1475;
 buffer[925] = 1474;
 buffer[926] = 1473;
 buffer[927] = 1472;
 buffer[928] = 1471;
 buffer[929] = 1470;
 buffer[930] = 1469;
 buffer[931] = 1468;
 buffer[932] = 1467;
 buffer[933] = 1466;
 buffer[934] = 1465;
 buffer[935] = 1464;
 buffer[936] = 1463;
 buffer[937] = 1462;
 buffer[938] = 1461;
 buffer[939] = 1460;
 buffer[940] = 1459;
 buffer[941] = 1458;
 buffer[942] = 1457;
 buffer[943] = 1456;
 buffer[944] = 1455;
 buffer[945] = 1454;
 buffer[946] = 1453;
 buffer[947] = 1452;
 buffer[948] = 1451;
 buffer[949] = 1450;
 buffer[950] = 1449;
 buffer[951] = 1448;
 buffer[952] = 1447;
 buffer[953] = 1446;
 buffer[954] = 1445;
 buffer[955] = 1444;
 buffer[956] = 1443;
 buffer[957] = 1442;
 buffer[958] = 1441;
 buffer[959] = 1440;
 buffer[960] = 1439;
 buffer[961] = 1438;
 buffer[962] = 1437;
 buffer[963] = 1436;
 buffer[964] = 1435;
 buffer[965] = 1434;
 buffer[966] = 1433;
 buffer[967] = 1432;
 buffer[968] = 1431;
 buffer[969] = 1430;
 buffer[970] = 1429;
 buffer[971] = 1428;
 buffer[972] = 1427;
 buffer[973] = 1426;
 buffer[974] = 1425;
 buffer[975] = 1424;
 buffer[976] = 1423;
 buffer[977] = 1422;
 buffer[978] = 1421;
 buffer[979] = 1420;
 buffer[980] = 1419;
 buffer[981] = 1418;
 buffer[982] = 1417;
 buffer[983] = 1416;
 buffer[984] = 1415;
 buffer[985] = 1414;
 buffer[986] = 1413;
 buffer[987] = 1412;
 buffer[988] = 1411;
 buffer[989] = 1410;
 buffer[990] = 1409;
 buffer[991] = 1408;
 buffer[992] = 1407;
 buffer[993] = 1406;
 buffer[994] = 1405;
 buffer[995] = 1404;
 buffer[996] = 1403;
 buffer[997] = 1402;
 buffer[998] = 1401;
 buffer[999] = 1400;
 buffer[1000] = 1399;
 buffer[1001] = 1398;
 buffer[1002] = 1397;
 buffer[1003] = 1396;
 buffer[1004] = 1395;
 buffer[1005] = 1394;
 buffer[1006] = 1393;
 buffer[1007] = 1392;
 buffer[1008] = 1391;
 buffer[1009] = 1390;
 buffer[1010] = 1389;
 buffer[1011] = 1388;
 buffer[1012] = 1387;
 buffer[1013] = 1386;
 buffer[1014] = 1385;
 buffer[1015] = 1384;
 buffer[1016] = 1383;
 buffer[1017] = 1382;
 buffer[1018] = 1381;
 buffer[1019] = 1380;
 buffer[1020] = 1379;
 buffer[1021] = 1378;
 buffer[1022] = 1377;
 buffer[1023] = 1376;
 buffer[1024] = 1375;
 buffer[1025] = 1374;
 buffer[1026] = 1373;
 buffer[1027] = 1372;
 buffer[1028] = 1371;
 buffer[1029] = 1370;
 buffer[1030] = 1369;
 buffer[1031] = 1368;
 buffer[1032] = 1367;
 buffer[1033] = 1366;
 buffer[1034] = 1365;
 buffer[1035] = 1364;
 buffer[1036] = 1363;
 buffer[1037] = 1362;
 buffer[1038] = 1361;
 buffer[1039] = 1360;
 buffer[1040] = 1359;
 buffer[1041] = 1358;
 buffer[1042] = 1357;
 buffer[1043] = 1356;
 buffer[1044] = 1355;
 buffer[1045] = 1354;
 buffer[1046] = 1353;
 buffer[1047] = 1352;
 buffer[1048] = 1351;
 buffer[1049] = 1350;
 buffer[1050] = 1349;
 buffer[1051] = 1348;
 buffer[1052] = 1347;
 buffer[1053] = 1346;
 buffer[1054] = 1345;
 buffer[1055] = 1344;
 buffer[1056] = 1343;
 buffer[1057] = 1342;
 buffer[1058] = 1341;
 buffer[1059] = 1340;
 buffer[1060] = 1339;
 buffer[1061] = 1338;
 buffer[1062] = 1337;
 buffer[1063] = 1336;
 buffer[1064] = 1335;
 buffer[1065] = 1334;
 buffer[1066] = 1333;
 buffer[1067] = 1332;
 buffer[1068] = 1331;
 buffer[1069] = 1330;
 buffer[1070] = 1329;
 buffer[1071] = 1328;
 buffer[1072] = 1327;
 buffer[1073] = 1326;
 buffer[1074] = 1325;
 buffer[1075] = 1324;
 buffer[1076] = 1323;
 buffer[1077] = 1322;
 buffer[1078] = 1321;
 buffer[1079] = 1320;
 buffer[1080] = 1319;
 buffer[1081] = 1318;
 buffer[1082] = 1317;
 buffer[1083] = 1316;
 buffer[1084] = 1315;
 buffer[1085] = 1314;
 buffer[1086] = 1313;
 buffer[1087] = 1312;
 buffer[1088] = 1311;
 buffer[1089] = 1310;
 buffer[1090] = 1309;
 buffer[1091] = 1308;
 buffer[1092] = 1307;
 buffer[1093] = 1306;
 buffer[1094] = 1305;
 buffer[1095] = 1304;
 buffer[1096] = 1303;
 buffer[1097] = 1302;
 buffer[1098] = 1301;
 buffer[1099] = 1300;
 buffer[1100] = 1299;
 buffer[1101] = 1298;
 buffer[1102] = 1297;
 buffer[1103] = 1296;
 buffer[1104] = 1295;
 buffer[1105] = 1294;
 buffer[1106] = 1293;
 buffer[1107] = 1292;
 buffer[1108] = 1291;
 buffer[1109] = 1290;
 buffer[1110] = 1289;
 buffer[1111] = 1288;
 buffer[1112] = 1287;
 buffer[1113] = 1286;
 buffer[1114] = 1285;
 buffer[1115] = 1284;
 buffer[1116] = 1283;
 buffer[1117] = 1282;
 buffer[1118] = 1281;
 buffer[1119] = 1280;
 buffer[1120] = 1279;
 buffer[1121] = 1278;
 buffer[1122] = 1277;
 buffer[1123] = 1276;
 buffer[1124] = 1275;
 buffer[1125] = 1274;
 buffer[1126] = 1273;
 buffer[1127] = 1272;
 buffer[1128] = 1271;
 buffer[1129] = 1270;
 buffer[1130] = 1269;
 buffer[1131] = 1268;
 buffer[1132] = 1267;
 buffer[1133] = 1266;
 buffer[1134] = 1265;
 buffer[1135] = 1264;
 buffer[1136] = 1263;
 buffer[1137] = 1262;
 buffer[1138] = 1261;
 buffer[1139] = 1260;
 buffer[1140] = 1259;
 buffer[1141] = 1258;
 buffer[1142] = 1257;
 buffer[1143] = 1256;
 buffer[1144] = 1255;
 buffer[1145] = 1254;
 buffer[1146] = 1253;
 buffer[1147] = 1252;
 buffer[1148] = 1251;
 buffer[1149] = 1250;
 buffer[1150] = 1249;
 buffer[1151] = 1248;
 buffer[1152] = 1247;
 buffer[1153] = 1246;
 buffer[1154] = 1245;
 buffer[1155] = 1244;
 buffer[1156] = 1243;
 buffer[1157] = 1242;
 buffer[1158] = 1241;
 buffer[1159] = 1240;
 buffer[1160] = 1239;
 buffer[1161] = 1238;
 buffer[1162] = 1237;
 buffer[1163] = 1236;
 buffer[1164] = 1235;
 buffer[1165] = 1234;
 buffer[1166] = 1233;
 buffer[1167] = 1232;
 buffer[1168] = 1231;
 buffer[1169] = 1230;
 buffer[1170] = 1229;
 buffer[1171] = 1228;
 buffer[1172] = 1227;
 buffer[1173] = 1226;
 buffer[1174] = 1225;
 buffer[1175] = 1224;
 buffer[1176] = 1223;
 buffer[1177] = 1222;
 buffer[1178] = 1221;
 buffer[1179] = 1220;
 buffer[1180] = 1219;
 buffer[1181] = 1218;
 buffer[1182] = 1217;
 buffer[1183] = 1216;
 buffer[1184] = 1215;
 buffer[1185] = 1214;
 buffer[1186] = 1213;
 buffer[1187] = 1212;
 buffer[1188] = 1211;
 buffer[1189] = 1210;
 buffer[1190] = 1209;
 buffer[1191] = 1208;
 buffer[1192] = 1207;
 buffer[1193] = 1206;
 buffer[1194] = 1205;
 buffer[1195] = 1204;
 buffer[1196] = 1203;
 buffer[1197] = 1202;
 buffer[1198] = 1201;
 buffer[1199] = 1200;
 buffer[1200] = 1199;
 buffer[1201] = 1198;
 buffer[1202] = 1197;
 buffer[1203] = 1196;
 buffer[1204] = 1195;
 buffer[1205] = 1194;
 buffer[1206] = 1193;
 buffer[1207] = 1192;
 buffer[1208] = 1191;
 buffer[1209] = 1190;
 buffer[1210] = 1189;
 buffer[1211] = 1188;
 buffer[1212] = 1187;
 buffer[1213] = 1186;
 buffer[1214] = 1185;
 buffer[1215] = 1184;
 buffer[1216] = 1183;
 buffer[1217] = 1182;
 buffer[1218] = 1181;
 buffer[1219] = 1180;
 buffer[1220] = 1179;
 buffer[1221] = 1178;
 buffer[1222] = 1177;
 buffer[1223] = 1176;
 buffer[1224] = 1175;
 buffer[1225] = 1174;
 buffer[1226] = 1173;
 buffer[1227] = 1172;
 buffer[1228] = 1171;
 buffer[1229] = 1170;
 buffer[1230] = 1169;
 buffer[1231] = 1168;
 buffer[1232] = 1167;
 buffer[1233] = 1166;
 buffer[1234] = 1165;
 buffer[1235] = 1164;
 buffer[1236] = 1163;
 buffer[1237] = 1162;
 buffer[1238] = 1161;
 buffer[1239] = 1160;
 buffer[1240] = 1159;
 buffer[1241] = 1158;
 buffer[1242] = 1157;
 buffer[1243] = 1156;
 buffer[1244] = 1155;
 buffer[1245] = 1154;
 buffer[1246] = 1153;
 buffer[1247] = 1152;
 buffer[1248] = 1151;
 buffer[1249] = 1150;
 buffer[1250] = 1149;
 buffer[1251] = 1148;
 buffer[1252] = 1147;
 buffer[1253] = 1146;
 buffer[1254] = 1145;
 buffer[1255] = 1144;
 buffer[1256] = 1143;
 buffer[1257] = 1142;
 buffer[1258] = 1141;
 buffer[1259] = 1140;
 buffer[1260] = 1139;
 buffer[1261] = 1138;
 buffer[1262] = 1137;
 buffer[1263] = 1136;
 buffer[1264] = 1135;
 buffer[1265] = 1134;
 buffer[1266] = 1133;
 buffer[1267] = 1132;
 buffer[1268] = 1131;
 buffer[1269] = 1130;
 buffer[1270] = 1129;
 buffer[1271] = 1128;
 buffer[1272] = 1127;
 buffer[1273] = 1126;
 buffer[1274] = 1125;
 buffer[1275] = 1124;
 buffer[1276] = 1123;
 buffer[1277] = 1122;
 buffer[1278] = 1121;
 buffer[1279] = 1120;
 buffer[1280] = 1119;
 buffer[1281] = 1118;
 buffer[1282] = 1117;
 buffer[1283] = 1116;
 buffer[1284] = 1115;
 buffer[1285] = 1114;
 buffer[1286] = 1113;
 buffer[1287] = 1112;
 buffer[1288] = 1111;
 buffer[1289] = 1110;
 buffer[1290] = 1109;
 buffer[1291] = 1108;
 buffer[1292] = 1107;
 buffer[1293] = 1106;
 buffer[1294] = 1105;
 buffer[1295] = 1104;
 buffer[1296] = 1103;
 buffer[1297] = 1102;
 buffer[1298] = 1101;
 buffer[1299] = 1100;
 buffer[1300] = 1099;
 buffer[1301] = 1098;
 buffer[1302] = 1097;
 buffer[1303] = 1096;
 buffer[1304] = 1095;
 buffer[1305] = 1094;
 buffer[1306] = 1093;
 buffer[1307] = 1092;
 buffer[1308] = 1091;
 buffer[1309] = 1090;
 buffer[1310] = 1089;
 buffer[1311] = 1088;
 buffer[1312] = 1087;
 buffer[1313] = 1086;
 buffer[1314] = 1085;
 buffer[1315] = 1084;
 buffer[1316] = 1083;
 buffer[1317] = 1082;
 buffer[1318] = 1081;
 buffer[1319] = 1080;
 buffer[1320] = 1079;
 buffer[1321] = 1078;
 buffer[1322] = 1077;
 buffer[1323] = 1076;
 buffer[1324] = 1075;
 buffer[1325] = 1074;
 buffer[1326] = 1073;
 buffer[1327] = 1072;
 buffer[1328] = 1071;
 buffer[1329] = 1070;
 buffer[1330] = 1069;
 buffer[1331] = 1068;
 buffer[1332] = 1067;
 buffer[1333] = 1066;
 buffer[1334] = 1065;
 buffer[1335] = 1064;
 buffer[1336] = 1063;
 buffer[1337] = 1062;
 buffer[1338] = 1061;
 buffer[1339] = 1060;
 buffer[1340] = 1059;
 buffer[1341] = 1058;
 buffer[1342] = 1057;
 buffer[1343] = 1056;
 buffer[1344] = 1055;
 buffer[1345] = 1054;
 buffer[1346] = 1053;
 buffer[1347] = 1052;
 buffer[1348] = 1051;
 buffer[1349] = 1050;
 buffer[1350] = 1049;
 buffer[1351] = 1048;
 buffer[1352] = 1047;
 buffer[1353] = 1046;
 buffer[1354] = 1045;
 buffer[1355] = 1044;
 buffer[1356] = 1043;
 buffer[1357] = 1042;
 buffer[1358] = 1041;
 buffer[1359] = 1040;
 buffer[1360] = 1039;
 buffer[1361] = 1038;
 buffer[1362] = 1037;
 buffer[1363] = 1036;
 buffer[1364] = 1035;
 buffer[1365] = 1034;
 buffer[1366] = 1033;
 buffer[1367] = 1032;
 buffer[1368] = 1031;
 buffer[1369] = 1030;
 buffer[1370] = 1029;
 buffer[1371] = 1028;
 buffer[1372] = 1027;
 buffer[1373] = 1026;
 buffer[1374] = 1025;
 buffer[1375] = 1024;
 buffer[1376] = 1023;
 buffer[1377] = 1022;
 buffer[1378] = 1021;
 buffer[1379] = 1020;
 buffer[1380] = 1019;
 buffer[1381] = 1018;
 buffer[1382] = 1017;
 buffer[1383] = 1016;
 buffer[1384] = 1015;
 buffer[1385] = 1014;
 buffer[1386] = 1013;
 buffer[1387] = 1012;
 buffer[1388] = 1011;
 buffer[1389] = 1010;
 buffer[1390] = 1009;
 buffer[1391] = 1008;
 buffer[1392] = 1007;
 buffer[1393] = 1006;
 buffer[1394] = 1005;
 buffer[1395] = 1004;
 buffer[1396] = 1003;
 buffer[1397] = 1002;
 buffer[1398] = 1001;
 buffer[1399] = 1000;
 buffer[1400] = 999;
 buffer[1401] = 998;
 buffer[1402] = 997;
 buffer[1403] = 996;
 buffer[1404] = 995;
 buffer[1405] = 994;
 buffer[1406] = 993;
 buffer[1407] = 992;
 buffer[1408] = 991;
 buffer[1409] = 990;
 buffer[1410] = 989;
 buffer[1411] = 988;
 buffer[1412] = 987;
 buffer[1413] = 986;
 buffer[1414] = 985;
 buffer[1415] = 984;
 buffer[1416] = 983;
 buffer[1417] = 982;
 buffer[1418] = 981;
 buffer[1419] = 980;
 buffer[1420] = 979;
 buffer[1421] = 978;
 buffer[1422] = 977;
 buffer[1423] = 976;
 buffer[1424] = 975;
 buffer[1425] = 974;
 buffer[1426] = 973;
 buffer[1427] = 972;
 buffer[1428] = 971;
 buffer[1429] = 970;
 buffer[1430] = 969;
 buffer[1431] = 968;
 buffer[1432] = 967;
 buffer[1433] = 966;
 buffer[1434] = 965;
 buffer[1435] = 964;
 buffer[1436] = 963;
 buffer[1437] = 962;
 buffer[1438] = 961;
 buffer[1439] = 960;
 buffer[1440] = 959;
 buffer[1441] = 958;
 buffer[1442] = 957;
 buffer[1443] = 956;
 buffer[1444] = 955;
 buffer[1445] = 954;
 buffer[1446] = 953;
 buffer[1447] = 952;
 buffer[1448] = 951;
 buffer[1449] = 950;
 buffer[1450] = 949;
 buffer[1451] = 948;
 buffer[1452] = 947;
 buffer[1453] = 946;
 buffer[1454] = 945;
 buffer[1455] = 944;
 buffer[1456] = 943;
 buffer[1457] = 942;
 buffer[1458] = 941;
 buffer[1459] = 940;
 buffer[1460] = 939;
 buffer[1461] = 938;
 buffer[1462] = 937;
 buffer[1463] = 936;
 buffer[1464] = 935;
 buffer[1465] = 934;
 buffer[1466] = 933;
 buffer[1467] = 932;
 buffer[1468] = 931;
 buffer[1469] = 930;
 buffer[1470] = 929;
 buffer[1471] = 928;
 buffer[1472] = 927;
 buffer[1473] = 926;
 buffer[1474] = 925;
 buffer[1475] = 924;
 buffer[1476] = 923;
 buffer[1477] = 922;
 buffer[1478] = 921;
 buffer[1479] = 920;
 buffer[1480] = 919;
 buffer[1481] = 918;
 buffer[1482] = 917;
 buffer[1483] = 916;
 buffer[1484] = 915;
 buffer[1485] = 914;
 buffer[1486] = 913;
 buffer[1487] = 912;
 buffer[1488] = 911;
 buffer[1489] = 910;
 buffer[1490] = 909;
 buffer[1491] = 908;
 buffer[1492] = 907;
 buffer[1493] = 906;
 buffer[1494] = 905;
 buffer[1495] = 904;
 buffer[1496] = 903;
 buffer[1497] = 902;
 buffer[1498] = 901;
 buffer[1499] = 900;
 buffer[1500] = 899;
 buffer[1501] = 898;
 buffer[1502] = 897;
 buffer[1503] = 896;
 buffer[1504] = 895;
 buffer[1505] = 894;
 buffer[1506] = 893;
 buffer[1507] = 892;
 buffer[1508] = 891;
 buffer[1509] = 890;
 buffer[1510] = 889;
 buffer[1511] = 888;
 buffer[1512] = 887;
 buffer[1513] = 886;
 buffer[1514] = 885;
 buffer[1515] = 884;
 buffer[1516] = 883;
 buffer[1517] = 882;
 buffer[1518] = 881;
 buffer[1519] = 880;
 buffer[1520] = 879;
 buffer[1521] = 878;
 buffer[1522] = 877;
 buffer[1523] = 876;
 buffer[1524] = 875;
 buffer[1525] = 874;
 buffer[1526] = 873;
 buffer[1527] = 872;
 buffer[1528] = 871;
 buffer[1529] = 870;
 buffer[1530] = 869;
 buffer[1531] = 868;
 buffer[1532] = 867;
 buffer[1533] = 866;
 buffer[1534] = 865;
 buffer[1535] = 864;
 buffer[1536] = 863;
 buffer[1537] = 862;
 buffer[1538] = 861;
 buffer[1539] = 860;
 buffer[1540] = 859;
 buffer[1541] = 858;
 buffer[1542] = 857;
 buffer[1543] = 856;
 buffer[1544] = 855;
 buffer[1545] = 854;
 buffer[1546] = 853;
 buffer[1547] = 852;
 buffer[1548] = 851;
 buffer[1549] = 850;
 buffer[1550] = 849;
 buffer[1551] = 848;
 buffer[1552] = 847;
 buffer[1553] = 846;
 buffer[1554] = 845;
 buffer[1555] = 844;
 buffer[1556] = 843;
 buffer[1557] = 842;
 buffer[1558] = 841;
 buffer[1559] = 840;
 buffer[1560] = 839;
 buffer[1561] = 838;
 buffer[1562] = 837;
 buffer[1563] = 836;
 buffer[1564] = 835;
 buffer[1565] = 834;
 buffer[1566] = 833;
 buffer[1567] = 832;
 buffer[1568] = 831;
 buffer[1569] = 830;
 buffer[1570] = 829;
 buffer[1571] = 828;
 buffer[1572] = 827;
 buffer[1573] = 826;
 buffer[1574] = 825;
 buffer[1575] = 824;
 buffer[1576] = 823;
 buffer[1577] = 822;
 buffer[1578] = 821;
 buffer[1579] = 820;
 buffer[1580] = 819;
 buffer[1581] = 818;
 buffer[1582] = 817;
 buffer[1583] = 816;
 buffer[1584] = 815;
 buffer[1585] = 814;
 buffer[1586] = 813;
 buffer[1587] = 812;
 buffer[1588] = 811;
 buffer[1589] = 810;
 buffer[1590] = 809;
 buffer[1591] = 808;
 buffer[1592] = 807;
 buffer[1593] = 806;
 buffer[1594] = 805;
 buffer[1595] = 804;
 buffer[1596] = 803;
 buffer[1597] = 802;
 buffer[1598] = 801;
 buffer[1599] = 800;
 buffer[1600] = 799;
 buffer[1601] = 798;
 buffer[1602] = 797;
 buffer[1603] = 796;
 buffer[1604] = 795;
 buffer[1605] = 794;
 buffer[1606] = 793;
 buffer[1607] = 792;
 buffer[1608] = 791;
 buffer[1609] = 790;
 buffer[1610] = 789;
 buffer[1611] = 788;
 buffer[1612] = 787;
 buffer[1613] = 786;
 buffer[1614] = 785;
 buffer[1615] = 784;
 buffer[1616] = 783;
 buffer[1617] = 782;
 buffer[1618] = 781;
 buffer[1619] = 780;
 buffer[1620] = 779;
 buffer[1621] = 778;
 buffer[1622] = 777;
 buffer[1623] = 776;
 buffer[1624] = 775;
 buffer[1625] = 774;
 buffer[1626] = 773;
 buffer[1627] = 772;
 buffer[1628] = 771;
 buffer[1629] = 770;
 buffer[1630] = 769;
 buffer[1631] = 768;
 buffer[1632] = 767;
 buffer[1633] = 766;
 buffer[1634] = 765;
 buffer[1635] = 764;
 buffer[1636] = 763;
 buffer[1637] = 762;
 buffer[1638] = 761;
 buffer[1639] = 760;
 buffer[1640] = 759;
 buffer[1641] = 758;
 buffer[1642] = 757;
 buffer[1643] = 756;
 buffer[1644] = 755;
 buffer[1645] = 754;
 buffer[1646] = 753;
 buffer[1647] = 752;
 buffer[1648] = 751;
 buffer[1649] = 750;
 buffer[1650] = 749;
 buffer[1651] = 748;
 buffer[1652] = 747;
 buffer[1653] = 746;
 buffer[1654] = 745;
 buffer[1655] = 744;
 buffer[1656] = 743;
 buffer[1657] = 742;
 buffer[1658] = 741;
 buffer[1659] = 740;
 buffer[1660] = 739;
 buffer[1661] = 738;
 buffer[1662] = 737;
 buffer[1663] = 736;
 buffer[1664] = 735;
 buffer[1665] = 734;
 buffer[1666] = 733;
 buffer[1667] = 732;
 buffer[1668] = 731;
 buffer[1669] = 730;
 buffer[1670] = 729;
 buffer[1671] = 728;
 buffer[1672] = 727;
 buffer[1673] = 726;
 buffer[1674] = 725;
 buffer[1675] = 724;
 buffer[1676] = 723;
 buffer[1677] = 722;
 buffer[1678] = 721;
 buffer[1679] = 720;
 buffer[1680] = 719;
 buffer[1681] = 718;
 buffer[1682] = 717;
 buffer[1683] = 716;
 buffer[1684] = 715;
 buffer[1685] = 714;
 buffer[1686] = 713;
 buffer[1687] = 712;
 buffer[1688] = 711;
 buffer[1689] = 710;
 buffer[1690] = 709;
 buffer[1691] = 708;
 buffer[1692] = 707;
 buffer[1693] = 706;
 buffer[1694] = 705;
 buffer[1695] = 704;
 buffer[1696] = 703;
 buffer[1697] = 702;
 buffer[1698] = 701;
 buffer[1699] = 700;
 buffer[1700] = 699;
 buffer[1701] = 698;
 buffer[1702] = 697;
 buffer[1703] = 696;
 buffer[1704] = 695;
 buffer[1705] = 694;
 buffer[1706] = 693;
 buffer[1707] = 692;
 buffer[1708] = 691;
 buffer[1709] = 690;
 buffer[1710] = 689;
 buffer[1711] = 688;
 buffer[1712] = 687;
 buffer[1713] = 686;
 buffer[1714] = 685;
 buffer[1715] = 684;
 buffer[1716] = 683;
 buffer[1717] = 682;
 buffer[1718] = 681;
 buffer[1719] = 680;
 buffer[1720] = 679;
 buffer[1721] = 678;
 buffer[1722] = 677;
 buffer[1723] = 676;
 buffer[1724] = 675;
 buffer[1725] = 674;
 buffer[1726] = 673;
 buffer[1727] = 672;
 buffer[1728] = 671;
 buffer[1729] = 670;
 buffer[1730] = 669;
 buffer[1731] = 668;
 buffer[1732] = 667;
 buffer[1733] = 666;
 buffer[1734] = 665;
 buffer[1735] = 664;
 buffer[1736] = 663;
 buffer[1737] = 662;
 buffer[1738] = 661;
 buffer[1739] = 660;
 buffer[1740] = 659;
 buffer[1741] = 658;
 buffer[1742] = 657;
 buffer[1743] = 656;
 buffer[1744] = 655;
 buffer[1745] = 654;
 buffer[1746] = 653;
 buffer[1747] = 652;
 buffer[1748] = 651;
 buffer[1749] = 650;
 buffer[1750] = 649;
 buffer[1751] = 648;
 buffer[1752] = 647;
 buffer[1753] = 646;
 buffer[1754] = 645;
 buffer[1755] = 644;
 buffer[1756] = 643;
 buffer[1757] = 642;
 buffer[1758] = 641;
 buffer[1759] = 640;
 buffer[1760] = 639;
 buffer[1761] = 638;
 buffer[1762] = 637;
 buffer[1763] = 636;
 buffer[1764] = 635;
 buffer[1765] = 634;
 buffer[1766] = 633;
 buffer[1767] = 632;
 buffer[1768] = 631;
 buffer[1769] = 630;
 buffer[1770] = 629;
 buffer[1771] = 628;
 buffer[1772] = 627;
 buffer[1773] = 626;
 buffer[1774] = 625;
 buffer[1775] = 624;
 buffer[1776] = 623;
 buffer[1777] = 622;
 buffer[1778] = 621;
 buffer[1779] = 620;
 buffer[1780] = 619;
 buffer[1781] = 618;
 buffer[1782] = 617;
 buffer[1783] = 616;
 buffer[1784] = 615;
 buffer[1785] = 614;
 buffer[1786] = 613;
 buffer[1787] = 612;
 buffer[1788] = 611;
 buffer[1789] = 610;
 buffer[1790] = 609;
 buffer[1791] = 608;
 buffer[1792] = 607;
 buffer[1793] = 606;
 buffer[1794] = 605;
 buffer[1795] = 604;
 buffer[1796] = 603;
 buffer[1797] = 602;
 buffer[1798] = 601;
 buffer[1799] = 600;
 buffer[1800] = 599;
 buffer[1801] = 598;
 buffer[1802] = 597;
 buffer[1803] = 596;
 buffer[1804] = 595;
 buffer[1805] = 594;
 buffer[1806] = 593;
 buffer[1807] = 592;
 buffer[1808] = 591;
 buffer[1809] = 590;
 buffer[1810] = 589;
 buffer[1811] = 588;
 buffer[1812] = 587;
 buffer[1813] = 586;
 buffer[1814] = 585;
 buffer[1815] = 584;
 buffer[1816] = 583;
 buffer[1817] = 582;
 buffer[1818] = 581;
 buffer[1819] = 580;
 buffer[1820] = 579;
 buffer[1821] = 578;
 buffer[1822] = 577;
 buffer[1823] = 576;
 buffer[1824] = 575;
 buffer[1825] = 574;
 buffer[1826] = 573;
 buffer[1827] = 572;
 buffer[1828] = 571;
 buffer[1829] = 570;
 buffer[1830] = 569;
 buffer[1831] = 568;
 buffer[1832] = 567;
 buffer[1833] = 566;
 buffer[1834] = 565;
 buffer[1835] = 564;
 buffer[1836] = 563;
 buffer[1837] = 562;
 buffer[1838] = 561;
 buffer[1839] = 560;
 buffer[1840] = 559;
 buffer[1841] = 558;
 buffer[1842] = 557;
 buffer[1843] = 556;
 buffer[1844] = 555;
 buffer[1845] = 554;
 buffer[1846] = 553;
 buffer[1847] = 552;
 buffer[1848] = 551;
 buffer[1849] = 550;
 buffer[1850] = 549;
 buffer[1851] = 548;
 buffer[1852] = 547;
 buffer[1853] = 546;
 buffer[1854] = 545;
 buffer[1855] = 544;
 buffer[1856] = 543;
 buffer[1857] = 542;
 buffer[1858] = 541;
 buffer[1859] = 540;
 buffer[1860] = 539;
 buffer[1861] = 538;
 buffer[1862] = 537;
 buffer[1863] = 536;
 buffer[1864] = 535;
 buffer[1865] = 534;
 buffer[1866] = 533;
 buffer[1867] = 532;
 buffer[1868] = 531;
 buffer[1869] = 530;
 buffer[1870] = 529;
 buffer[1871] = 528;
 buffer[1872] = 527;
 buffer[1873] = 526;
 buffer[1874] = 525;
 buffer[1875] = 524;
 buffer[1876] = 523;
 buffer[1877] = 522;
 buffer[1878] = 521;
 buffer[1879] = 520;
 buffer[1880] = 519;
 buffer[1881] = 518;
 buffer[1882] = 517;
 buffer[1883] = 516;
 buffer[1884] = 515;
 buffer[1885] = 514;
 buffer[1886] = 513;
 buffer[1887] = 512;
 buffer[1888] = 511;
 buffer[1889] = 510;
 buffer[1890] = 509;
 buffer[1891] = 508;
 buffer[1892] = 507;
 buffer[1893] = 506;
 buffer[1894] = 505;
 buffer[1895] = 504;
 buffer[1896] = 503;
 buffer[1897] = 502;
 buffer[1898] = 501;
 buffer[1899] = 500;
 buffer[1900] = 499;
 buffer[1901] = 498;
 buffer[1902] = 497;
 buffer[1903] = 496;
 buffer[1904] = 495;
 buffer[1905] = 494;
 buffer[1906] = 493;
 buffer[1907] = 492;
 buffer[1908] = 491;
 buffer[1909] = 490;
 buffer[1910] = 489;
 buffer[1911] = 488;
 buffer[1912] = 487;
 buffer[1913] = 486;
 buffer[1914] = 485;
 buffer[1915] = 484;
 buffer[1916] = 483;
 buffer[1917] = 482;
 buffer[1918] = 481;
 buffer[1919] = 480;
 buffer[1920] = 479;
 buffer[1921] = 478;
 buffer[1922] = 477;
 buffer[1923] = 476;
 buffer[1924] = 475;
 buffer[1925] = 474;
 buffer[1926] = 473;
 buffer[1927] = 472;
 buffer[1928] = 471;
 buffer[1929] = 470;
 buffer[1930] = 469;
 buffer[1931] = 468;
 buffer[1932] = 467;
 buffer[1933] = 466;
 buffer[1934] = 465;
 buffer[1935] = 464;
 buffer[1936] = 463;
 buffer[1937] = 462;
 buffer[1938] = 461;
 buffer[1939] = 460;
 buffer[1940] = 459;
 buffer[1941] = 458;
 buffer[1942] = 457;
 buffer[1943] = 456;
 buffer[1944] = 455;
 buffer[1945] = 454;
 buffer[1946] = 453;
 buffer[1947] = 452;
 buffer[1948] = 451;
 buffer[1949] = 450;
 buffer[1950] = 449;
 buffer[1951] = 448;
 buffer[1952] = 447;
 buffer[1953] = 446;
 buffer[1954] = 445;
 buffer[1955] = 444;
 buffer[1956] = 443;
 buffer[1957] = 442;
 buffer[1958] = 441;
 buffer[1959] = 440;
 buffer[1960] = 439;
 buffer[1961] = 438;
 buffer[1962] = 437;
 buffer[1963] = 436;
 buffer[1964] = 435;
 buffer[1965] = 434;
 buffer[1966] = 433;
 buffer[1967] = 432;
 buffer[1968] = 431;
 buffer[1969] = 430;
 buffer[1970] = 429;
 buffer[1971] = 428;
 buffer[1972] = 427;
 buffer[1973] = 426;
 buffer[1974] = 425;
 buffer[1975] = 424;
 buffer[1976] = 423;
 buffer[1977] = 422;
 buffer[1978] = 421;
 buffer[1979] = 420;
 buffer[1980] = 419;
 buffer[1981] = 418;
 buffer[1982] = 417;
 buffer[1983] = 416;
 buffer[1984] = 415;
 buffer[1985] = 414;
 buffer[1986] = 413;
 buffer[1987] = 412;
 buffer[1988] = 411;
 buffer[1989] = 410;
 buffer[1990] = 409;
 buffer[1991] = 408;
 buffer[1992] = 407;
 buffer[1993] = 406;
 buffer[1994] = 405;
 buffer[1995] = 404;
 buffer[1996] = 403;
 buffer[1997] = 402;
 buffer[1998] = 401;
 buffer[1999] = 400;
 buffer[2000] = 399;
 buffer[2001] = 398;
 buffer[2002] = 397;
 buffer[2003] = 396;
 buffer[2004] = 395;
 buffer[2005] = 394;
 buffer[2006] = 393;
 buffer[2007] = 392;
 buffer[2008] = 391;
 buffer[2009] = 390;
 buffer[2010] = 389;
 buffer[2011] = 388;
 buffer[2012] = 387;
 buffer[2013] = 386;
 buffer[2014] = 385;
 buffer[2015] = 384;
 buffer[2016] = 383;
 buffer[2017] = 382;
 buffer[2018] = 381;
 buffer[2019] = 380;
 buffer[2020] = 379;
 buffer[2021] = 378;
 buffer[2022] = 377;
 buffer[2023] = 376;
 buffer[2024] = 375;
 buffer[2025] = 374;
 buffer[2026] = 373;
 buffer[2027] = 372;
 buffer[2028] = 371;
 buffer[2029] = 370;
 buffer[2030] = 369;
 buffer[2031] = 368;
 buffer[2032] = 367;
 buffer[2033] = 366;
 buffer[2034] = 365;
 buffer[2035] = 364;
 buffer[2036] = 363;
 buffer[2037] = 362;
 buffer[2038] = 361;
 buffer[2039] = 360;
 buffer[2040] = 359;
 buffer[2041] = 358;
 buffer[2042] = 357;
 buffer[2043] = 356;
 buffer[2044] = 355;
 buffer[2045] = 354;
 buffer[2046] = 353;
 buffer[2047] = 352;
 buffer[2048] = 351;
 buffer[2049] = 350;
 buffer[2050] = 349;
 buffer[2051] = 348;
 buffer[2052] = 347;
 buffer[2053] = 346;
 buffer[2054] = 345;
 buffer[2055] = 344;
 buffer[2056] = 343;
 buffer[2057] = 342;
 buffer[2058] = 341;
 buffer[2059] = 340;
 buffer[2060] = 339;
 buffer[2061] = 338;
 buffer[2062] = 337;
 buffer[2063] = 336;
 buffer[2064] = 335;
 buffer[2065] = 334;
 buffer[2066] = 333;
 buffer[2067] = 332;
 buffer[2068] = 331;
 buffer[2069] = 330;
 buffer[2070] = 329;
 buffer[2071] = 328;
 buffer[2072] = 327;
 buffer[2073] = 326;
 buffer[2074] = 325;
 buffer[2075] = 324;
 buffer[2076] = 323;
 buffer[2077] = 322;
 buffer[2078] = 321;
 buffer[2079] = 320;
 buffer[2080] = 319;
 buffer[2081] = 318;
 buffer[2082] = 317;
 buffer[2083] = 316;
 buffer[2084] = 315;
 buffer[2085] = 314;
 buffer[2086] = 313;
 buffer[2087] = 312;
 buffer[2088] = 311;
 buffer[2089] = 310;
 buffer[2090] = 309;
 buffer[2091] = 308;
 buffer[2092] = 307;
 buffer[2093] = 306;
 buffer[2094] = 305;
 buffer[2095] = 304;
 buffer[2096] = 303;
 buffer[2097] = 302;
 buffer[2098] = 301;
 buffer[2099] = 300;
 buffer[2100] = 299;
 buffer[2101] = 298;
 buffer[2102] = 297;
 buffer[2103] = 296;
 buffer[2104] = 295;
 buffer[2105] = 294;
 buffer[2106] = 293;
 buffer[2107] = 292;
 buffer[2108] = 291;
 buffer[2109] = 290;
 buffer[2110] = 289;
 buffer[2111] = 288;
 buffer[2112] = 287;
 buffer[2113] = 286;
 buffer[2114] = 285;
 buffer[2115] = 284;
 buffer[2116] = 283;
 buffer[2117] = 282;
 buffer[2118] = 281;
 buffer[2119] = 280;
 buffer[2120] = 279;
 buffer[2121] = 278;
 buffer[2122] = 277;
 buffer[2123] = 276;
 buffer[2124] = 275;
 buffer[2125] = 274;
 buffer[2126] = 273;
 buffer[2127] = 272;
 buffer[2128] = 271;
 buffer[2129] = 270;
 buffer[2130] = 269;
 buffer[2131] = 268;
 buffer[2132] = 267;
 buffer[2133] = 266;
 buffer[2134] = 265;
 buffer[2135] = 264;
 buffer[2136] = 263;
 buffer[2137] = 262;
 buffer[2138] = 261;
 buffer[2139] = 260;
 buffer[2140] = 259;
 buffer[2141] = 258;
 buffer[2142] = 257;
 buffer[2143] = 256;
 buffer[2144] = 255;
 buffer[2145] = 254;
 buffer[2146] = 253;
 buffer[2147] = 252;
 buffer[2148] = 251;
 buffer[2149] = 250;
 buffer[2150] = 249;
 buffer[2151] = 248;
 buffer[2152] = 247;
 buffer[2153] = 246;
 buffer[2154] = 245;
 buffer[2155] = 244;
 buffer[2156] = 243;
 buffer[2157] = 242;
 buffer[2158] = 241;
 buffer[2159] = 240;
 buffer[2160] = 239;
 buffer[2161] = 238;
 buffer[2162] = 237;
 buffer[2163] = 236;
 buffer[2164] = 235;
 buffer[2165] = 234;
 buffer[2166] = 233;
 buffer[2167] = 232;
 buffer[2168] = 231;
 buffer[2169] = 230;
 buffer[2170] = 229;
 buffer[2171] = 228;
 buffer[2172] = 227;
 buffer[2173] = 226;
 buffer[2174] = 225;
 buffer[2175] = 224;
 buffer[2176] = 223;
 buffer[2177] = 222;
 buffer[2178] = 221;
 buffer[2179] = 220;
 buffer[2180] = 219;
 buffer[2181] = 218;
 buffer[2182] = 217;
 buffer[2183] = 216;
 buffer[2184] = 215;
 buffer[2185] = 214;
 buffer[2186] = 213;
 buffer[2187] = 212;
 buffer[2188] = 211;
 buffer[2189] = 210;
 buffer[2190] = 209;
 buffer[2191] = 208;
 buffer[2192] = 207;
 buffer[2193] = 206;
 buffer[2194] = 205;
 buffer[2195] = 204;
 buffer[2196] = 203;
 buffer[2197] = 202;
 buffer[2198] = 201;
 buffer[2199] = 200;
 buffer[2200] = 199;
 buffer[2201] = 198;
 buffer[2202] = 197;
 buffer[2203] = 196;
 buffer[2204] = 195;
 buffer[2205] = 194;
 buffer[2206] = 193;
 buffer[2207] = 192;
 buffer[2208] = 191;
 buffer[2209] = 190;
 buffer[2210] = 189;
 buffer[2211] = 188;
 buffer[2212] = 187;
 buffer[2213] = 186;
 buffer[2214] = 185;
 buffer[2215] = 184;
 buffer[2216] = 183;
 buffer[2217] = 182;
 buffer[2218] = 181;
 buffer[2219] = 180;
 buffer[2220] = 179;
 buffer[2221] = 178;
 buffer[2222] = 177;
 buffer[2223] = 176;
 buffer[2224] = 175;
 buffer[2225] = 174;
 buffer[2226] = 173;
 buffer[2227] = 172;
 buffer[2228] = 171;
 buffer[2229] = 170;
 buffer[2230] = 169;
 buffer[2231] = 168;
 buffer[2232] = 167;
 buffer[2233] = 166;
 buffer[2234] = 165;
 buffer[2235] = 164;
 buffer[2236] = 163;
 buffer[2237] = 162;
 buffer[2238] = 161;
 buffer[2239] = 160;
 buffer[2240] = 159;
 buffer[2241] = 158;
 buffer[2242] = 157;
 buffer[2243] = 156;
 buffer[2244] = 155;
 buffer[2245] = 154;
 buffer[2246] = 153;
 buffer[2247] = 152;
 buffer[2248] = 151;
 buffer[2249] = 150;
 buffer[2250] = 149;
 buffer[2251] = 148;
 buffer[2252] = 147;
 buffer[2253] = 146;
 buffer[2254] = 145;
 buffer[2255] = 144;
 buffer[2256] = 143;
 buffer[2257] = 142;
 buffer[2258] = 141;
 buffer[2259] = 140;
 buffer[2260] = 139;
 buffer[2261] = 138;
 buffer[2262] = 137;
 buffer[2263] = 136;
 buffer[2264] = 135;
 buffer[2265] = 134;
 buffer[2266] = 133;
 buffer[2267] = 132;
 buffer[2268] = 131;
 buffer[2269] = 130;
 buffer[2270] = 129;
 buffer[2271] = 128;
 buffer[2272] = 127;
 buffer[2273] = 126;
 buffer[2274] = 125;
 buffer[2275] = 124;
 buffer[2276] = 123;
 buffer[2277] = 122;
 buffer[2278] = 121;
 buffer[2279] = 120;
 buffer[2280] = 119;
 buffer[2281] = 118;
 buffer[2282] = 117;
 buffer[2283] = 116;
 buffer[2284] = 115;
 buffer[2285] = 114;
 buffer[2286] = 113;
 buffer[2287] = 112;
 buffer[2288] = 111;
 buffer[2289] = 110;
 buffer[2290] = 109;
 buffer[2291] = 108;
 buffer[2292] = 107;
 buffer[2293] = 106;
 buffer[2294] = 105;
 buffer[2295] = 104;
 buffer[2296] = 103;
 buffer[2297] = 102;
 buffer[2298] = 101;
 buffer[2299] = 100;
 buffer[2300] = 99;
 buffer[2301] = 98;
 buffer[2302] = 97;
 buffer[2303] = 96;
 buffer[2304] = 95;
 buffer[2305] = 94;
 buffer[2306] = 93;
 buffer[2307] = 92;
 buffer[2308] = 91;
 buffer[2309] = 90;
 buffer[2310] = 89;
 buffer[2311] = 88;
 buffer[2312] = 87;
 buffer[2313] = 86;
 buffer[2314] = 85;
 buffer[2315] = 84;
 buffer[2316] = 83;
 buffer[2317] = 82;
 buffer[2318] = 81;
 buffer[2319] = 80;
 buffer[2320] = 79;
 buffer[2321] = 78;
 buffer[2322] = 77;
 buffer[2323] = 76;
 buffer[2324] = 75;
 buffer[2325] = 74;
 buffer[2326] = 73;
 buffer[2327] = 72;
 buffer[2328] = 71;
 buffer[2329] = 70;
 buffer[2330] = 69;
 buffer[2331] = 68;
 buffer[2332] = 67;
 buffer[2333] = 66;
 buffer[2334] = 65;
 buffer[2335] = 64;
 buffer[2336] = 63;
 buffer[2337] = 62;
 buffer[2338] = 61;
 buffer[2339] = 60;
 buffer[2340] = 59;
 buffer[2341] = 58;
 buffer[2342] = 57;
 buffer[2343] = 56;
 buffer[2344] = 55;
 buffer[2345] = 54;
 buffer[2346] = 53;
 buffer[2347] = 52;
 buffer[2348] = 51;
 buffer[2349] = 50;
 buffer[2350] = 49;
 buffer[2351] = 48;
 buffer[2352] = 47;
 buffer[2353] = 46;
 buffer[2354] = 45;
 buffer[2355] = 44;
 buffer[2356] = 43;
 buffer[2357] = 42;
 buffer[2358] = 41;
 buffer[2359] = 40;
 buffer[2360] = 39;
 buffer[2361] = 38;
 buffer[2362] = 37;
 buffer[2363] = 36;
 buffer[2364] = 35;
 buffer[2365] = 34;
 buffer[2366] = 33;
 buffer[2367] = 32;
 buffer[2368] = 31;
 buffer[2369] = 30;
 buffer[2370] = 29;
 buffer[2371] = 28;
 buffer[2372] = 27;
 buffer[2373] = 26;
 buffer[2374] = 25;
 buffer[2375] = 24;
 buffer[2376] = 23;
 buffer[2377] = 22;
 buffer[2378] = 21;
 buffer[2379] = 20;
 buffer[2380] = 19;
 buffer[2381] = 18;
 buffer[2382] = 17;
 buffer[2383] = 16;
 buffer[2384] = 15;
 buffer[2385] = 14;
 buffer[2386] = 13;
 buffer[2387] = 12;
 buffer[2388] = 11;
 buffer[2389] = 10;
 buffer[2390] = 9;
 buffer[2391] = 8;
 buffer[2392] = 7;
 buffer[2393] = 6;
 buffer[2394] = 5;
 buffer[2395] = 4;
 buffer[2396] = 3;
 buffer[2397] = 2;
 buffer[2398] = 1;
 buffer[2399] = 0;
end

endmodule

module M_multiplex_display_mem_bitmap(
input      [0:0]             in_bitmap_wenable0,
input       [7:0]     in_bitmap_wdata0,
input      [18:0]                in_bitmap_addr0,
input      [0:0]             in_bitmap_wenable1,
input      [7:0]                 in_bitmap_wdata1,
input      [18:0]                in_bitmap_addr1,
output reg  [7:0]     out_bitmap_rdata0,
output reg  [7:0]     out_bitmap_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[307199:0];
always @(posedge clock0) begin
  if (in_bitmap_wenable0) begin
    buffer[in_bitmap_addr0] <= in_bitmap_wdata0;
  end else begin
    out_bitmap_rdata0 <= buffer[in_bitmap_addr0];
  end
end
always @(posedge clock1) begin
  if (in_bitmap_wenable1) begin
    buffer[in_bitmap_addr1] <= in_bitmap_wdata1;
  end else begin
    out_bitmap_rdata1 <= buffer[in_bitmap_addr1];
  end
end

endmodule

module M_multiplex_display (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_gpu_x,
in_gpu_y,
in_gpu_dotset,
in_gpu_write,
in_tpu_x,
in_tpu_y,
in_tpu_set,
in_tpu_write,
out_pix_red,
out_pix_green,
out_pix_blue,
in_run,
out_done,
reset,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [9:0] in_gpu_x;
input  [8:0] in_gpu_y;
input  [7:0] in_gpu_dotset;
input  [0:0] in_gpu_write;
input  [6:0] in_tpu_x;
input  [4:0] in_tpu_y;
input  [7:0] in_tpu_set;
input  [1:0] in_tpu_write;
output  [5:0] out_pix_red;
output  [5:0] out_pix_green;
output  [5:0] out_pix_blue;
input in_run;
output out_done;
input reset;
input clock;
wire  [7:0] _w_mem_character_rdata0;
wire  [7:0] _w_mem_character_rdata1;
wire  [7:0] _w_mem_foreground_rdata0;
wire  [7:0] _w_mem_foreground_rdata1;
wire  [7:0] _w_mem_background_rdata0;
wire  [7:0] _w_mem_background_rdata1;
wire  [7:0] _w_mem_bitmap_rdata0;
wire  [7:0] _w_mem_bitmap_rdata1;
wire  [7:0] _c_characterGenerator[4095:0];
assign _c_characterGenerator[0] = 8'h00;
assign _c_characterGenerator[1] = 8'h00;
assign _c_characterGenerator[2] = 8'h00;
assign _c_characterGenerator[3] = 8'h00;
assign _c_characterGenerator[4] = 8'h00;
assign _c_characterGenerator[5] = 8'h00;
assign _c_characterGenerator[6] = 8'h00;
assign _c_characterGenerator[7] = 8'h00;
assign _c_characterGenerator[8] = 8'h00;
assign _c_characterGenerator[9] = 8'h00;
assign _c_characterGenerator[10] = 8'h00;
assign _c_characterGenerator[11] = 8'h00;
assign _c_characterGenerator[12] = 8'h00;
assign _c_characterGenerator[13] = 8'h00;
assign _c_characterGenerator[14] = 8'h00;
assign _c_characterGenerator[15] = 8'h00;
assign _c_characterGenerator[16] = 8'h00;
assign _c_characterGenerator[17] = 8'h00;
assign _c_characterGenerator[18] = 8'h7e;
assign _c_characterGenerator[19] = 8'h81;
assign _c_characterGenerator[20] = 8'ha5;
assign _c_characterGenerator[21] = 8'h81;
assign _c_characterGenerator[22] = 8'h81;
assign _c_characterGenerator[23] = 8'hbd;
assign _c_characterGenerator[24] = 8'h99;
assign _c_characterGenerator[25] = 8'h81;
assign _c_characterGenerator[26] = 8'h81;
assign _c_characterGenerator[27] = 8'h7e;
assign _c_characterGenerator[28] = 8'h00;
assign _c_characterGenerator[29] = 8'h00;
assign _c_characterGenerator[30] = 8'h00;
assign _c_characterGenerator[31] = 8'h00;
assign _c_characterGenerator[32] = 8'h00;
assign _c_characterGenerator[33] = 8'h00;
assign _c_characterGenerator[34] = 8'h7e;
assign _c_characterGenerator[35] = 8'hff;
assign _c_characterGenerator[36] = 8'hdb;
assign _c_characterGenerator[37] = 8'hff;
assign _c_characterGenerator[38] = 8'hff;
assign _c_characterGenerator[39] = 8'hc3;
assign _c_characterGenerator[40] = 8'he7;
assign _c_characterGenerator[41] = 8'hff;
assign _c_characterGenerator[42] = 8'hff;
assign _c_characterGenerator[43] = 8'h7e;
assign _c_characterGenerator[44] = 8'h00;
assign _c_characterGenerator[45] = 8'h00;
assign _c_characterGenerator[46] = 8'h00;
assign _c_characterGenerator[47] = 8'h00;
assign _c_characterGenerator[48] = 8'h00;
assign _c_characterGenerator[49] = 8'h00;
assign _c_characterGenerator[50] = 8'h00;
assign _c_characterGenerator[51] = 8'h00;
assign _c_characterGenerator[52] = 8'h6c;
assign _c_characterGenerator[53] = 8'hfe;
assign _c_characterGenerator[54] = 8'hfe;
assign _c_characterGenerator[55] = 8'hfe;
assign _c_characterGenerator[56] = 8'hfe;
assign _c_characterGenerator[57] = 8'h7c;
assign _c_characterGenerator[58] = 8'h38;
assign _c_characterGenerator[59] = 8'h10;
assign _c_characterGenerator[60] = 8'h00;
assign _c_characterGenerator[61] = 8'h00;
assign _c_characterGenerator[62] = 8'h00;
assign _c_characterGenerator[63] = 8'h00;
assign _c_characterGenerator[64] = 8'h00;
assign _c_characterGenerator[65] = 8'h00;
assign _c_characterGenerator[66] = 8'h00;
assign _c_characterGenerator[67] = 8'h00;
assign _c_characterGenerator[68] = 8'h10;
assign _c_characterGenerator[69] = 8'h38;
assign _c_characterGenerator[70] = 8'h7c;
assign _c_characterGenerator[71] = 8'hfe;
assign _c_characterGenerator[72] = 8'h7c;
assign _c_characterGenerator[73] = 8'h38;
assign _c_characterGenerator[74] = 8'h10;
assign _c_characterGenerator[75] = 8'h00;
assign _c_characterGenerator[76] = 8'h00;
assign _c_characterGenerator[77] = 8'h00;
assign _c_characterGenerator[78] = 8'h00;
assign _c_characterGenerator[79] = 8'h00;
assign _c_characterGenerator[80] = 8'h00;
assign _c_characterGenerator[81] = 8'h00;
assign _c_characterGenerator[82] = 8'h00;
assign _c_characterGenerator[83] = 8'h18;
assign _c_characterGenerator[84] = 8'h3c;
assign _c_characterGenerator[85] = 8'h3c;
assign _c_characterGenerator[86] = 8'he7;
assign _c_characterGenerator[87] = 8'he7;
assign _c_characterGenerator[88] = 8'he7;
assign _c_characterGenerator[89] = 8'h18;
assign _c_characterGenerator[90] = 8'h18;
assign _c_characterGenerator[91] = 8'h3c;
assign _c_characterGenerator[92] = 8'h00;
assign _c_characterGenerator[93] = 8'h00;
assign _c_characterGenerator[94] = 8'h00;
assign _c_characterGenerator[95] = 8'h00;
assign _c_characterGenerator[96] = 8'h00;
assign _c_characterGenerator[97] = 8'h00;
assign _c_characterGenerator[98] = 8'h00;
assign _c_characterGenerator[99] = 8'h18;
assign _c_characterGenerator[100] = 8'h3c;
assign _c_characterGenerator[101] = 8'h7e;
assign _c_characterGenerator[102] = 8'hff;
assign _c_characterGenerator[103] = 8'hff;
assign _c_characterGenerator[104] = 8'h7e;
assign _c_characterGenerator[105] = 8'h18;
assign _c_characterGenerator[106] = 8'h18;
assign _c_characterGenerator[107] = 8'h3c;
assign _c_characterGenerator[108] = 8'h00;
assign _c_characterGenerator[109] = 8'h00;
assign _c_characterGenerator[110] = 8'h00;
assign _c_characterGenerator[111] = 8'h00;
assign _c_characterGenerator[112] = 8'h00;
assign _c_characterGenerator[113] = 8'h00;
assign _c_characterGenerator[114] = 8'h00;
assign _c_characterGenerator[115] = 8'h00;
assign _c_characterGenerator[116] = 8'h00;
assign _c_characterGenerator[117] = 8'h00;
assign _c_characterGenerator[118] = 8'h18;
assign _c_characterGenerator[119] = 8'h3c;
assign _c_characterGenerator[120] = 8'h3c;
assign _c_characterGenerator[121] = 8'h18;
assign _c_characterGenerator[122] = 8'h00;
assign _c_characterGenerator[123] = 8'h00;
assign _c_characterGenerator[124] = 8'h00;
assign _c_characterGenerator[125] = 8'h00;
assign _c_characterGenerator[126] = 8'h00;
assign _c_characterGenerator[127] = 8'h00;
assign _c_characterGenerator[128] = 8'hff;
assign _c_characterGenerator[129] = 8'hff;
assign _c_characterGenerator[130] = 8'hff;
assign _c_characterGenerator[131] = 8'hff;
assign _c_characterGenerator[132] = 8'hff;
assign _c_characterGenerator[133] = 8'hff;
assign _c_characterGenerator[134] = 8'he7;
assign _c_characterGenerator[135] = 8'hc3;
assign _c_characterGenerator[136] = 8'hc3;
assign _c_characterGenerator[137] = 8'he7;
assign _c_characterGenerator[138] = 8'hff;
assign _c_characterGenerator[139] = 8'hff;
assign _c_characterGenerator[140] = 8'hff;
assign _c_characterGenerator[141] = 8'hff;
assign _c_characterGenerator[142] = 8'hff;
assign _c_characterGenerator[143] = 8'hff;
assign _c_characterGenerator[144] = 8'h00;
assign _c_characterGenerator[145] = 8'h00;
assign _c_characterGenerator[146] = 8'h00;
assign _c_characterGenerator[147] = 8'h00;
assign _c_characterGenerator[148] = 8'h00;
assign _c_characterGenerator[149] = 8'h3c;
assign _c_characterGenerator[150] = 8'h66;
assign _c_characterGenerator[151] = 8'h42;
assign _c_characterGenerator[152] = 8'h42;
assign _c_characterGenerator[153] = 8'h66;
assign _c_characterGenerator[154] = 8'h3c;
assign _c_characterGenerator[155] = 8'h00;
assign _c_characterGenerator[156] = 8'h00;
assign _c_characterGenerator[157] = 8'h00;
assign _c_characterGenerator[158] = 8'h00;
assign _c_characterGenerator[159] = 8'h00;
assign _c_characterGenerator[160] = 8'hff;
assign _c_characterGenerator[161] = 8'hff;
assign _c_characterGenerator[162] = 8'hff;
assign _c_characterGenerator[163] = 8'hff;
assign _c_characterGenerator[164] = 8'hff;
assign _c_characterGenerator[165] = 8'hc3;
assign _c_characterGenerator[166] = 8'h99;
assign _c_characterGenerator[167] = 8'hbd;
assign _c_characterGenerator[168] = 8'hbd;
assign _c_characterGenerator[169] = 8'h99;
assign _c_characterGenerator[170] = 8'hc3;
assign _c_characterGenerator[171] = 8'hff;
assign _c_characterGenerator[172] = 8'hff;
assign _c_characterGenerator[173] = 8'hff;
assign _c_characterGenerator[174] = 8'hff;
assign _c_characterGenerator[175] = 8'hff;
assign _c_characterGenerator[176] = 8'h00;
assign _c_characterGenerator[177] = 8'h00;
assign _c_characterGenerator[178] = 8'h1e;
assign _c_characterGenerator[179] = 8'h0e;
assign _c_characterGenerator[180] = 8'h1a;
assign _c_characterGenerator[181] = 8'h32;
assign _c_characterGenerator[182] = 8'h78;
assign _c_characterGenerator[183] = 8'hcc;
assign _c_characterGenerator[184] = 8'hcc;
assign _c_characterGenerator[185] = 8'hcc;
assign _c_characterGenerator[186] = 8'hcc;
assign _c_characterGenerator[187] = 8'h78;
assign _c_characterGenerator[188] = 8'h00;
assign _c_characterGenerator[189] = 8'h00;
assign _c_characterGenerator[190] = 8'h00;
assign _c_characterGenerator[191] = 8'h00;
assign _c_characterGenerator[192] = 8'h00;
assign _c_characterGenerator[193] = 8'h00;
assign _c_characterGenerator[194] = 8'h3c;
assign _c_characterGenerator[195] = 8'h66;
assign _c_characterGenerator[196] = 8'h66;
assign _c_characterGenerator[197] = 8'h66;
assign _c_characterGenerator[198] = 8'h66;
assign _c_characterGenerator[199] = 8'h3c;
assign _c_characterGenerator[200] = 8'h18;
assign _c_characterGenerator[201] = 8'h7e;
assign _c_characterGenerator[202] = 8'h18;
assign _c_characterGenerator[203] = 8'h18;
assign _c_characterGenerator[204] = 8'h00;
assign _c_characterGenerator[205] = 8'h00;
assign _c_characterGenerator[206] = 8'h00;
assign _c_characterGenerator[207] = 8'h00;
assign _c_characterGenerator[208] = 8'h00;
assign _c_characterGenerator[209] = 8'h00;
assign _c_characterGenerator[210] = 8'h3f;
assign _c_characterGenerator[211] = 8'h33;
assign _c_characterGenerator[212] = 8'h3f;
assign _c_characterGenerator[213] = 8'h30;
assign _c_characterGenerator[214] = 8'h30;
assign _c_characterGenerator[215] = 8'h30;
assign _c_characterGenerator[216] = 8'h30;
assign _c_characterGenerator[217] = 8'h70;
assign _c_characterGenerator[218] = 8'hf0;
assign _c_characterGenerator[219] = 8'he0;
assign _c_characterGenerator[220] = 8'h00;
assign _c_characterGenerator[221] = 8'h00;
assign _c_characterGenerator[222] = 8'h00;
assign _c_characterGenerator[223] = 8'h00;
assign _c_characterGenerator[224] = 8'h00;
assign _c_characterGenerator[225] = 8'h00;
assign _c_characterGenerator[226] = 8'h7f;
assign _c_characterGenerator[227] = 8'h63;
assign _c_characterGenerator[228] = 8'h7f;
assign _c_characterGenerator[229] = 8'h63;
assign _c_characterGenerator[230] = 8'h63;
assign _c_characterGenerator[231] = 8'h63;
assign _c_characterGenerator[232] = 8'h63;
assign _c_characterGenerator[233] = 8'h67;
assign _c_characterGenerator[234] = 8'he7;
assign _c_characterGenerator[235] = 8'he6;
assign _c_characterGenerator[236] = 8'hc0;
assign _c_characterGenerator[237] = 8'h00;
assign _c_characterGenerator[238] = 8'h00;
assign _c_characterGenerator[239] = 8'h00;
assign _c_characterGenerator[240] = 8'h00;
assign _c_characterGenerator[241] = 8'h00;
assign _c_characterGenerator[242] = 8'h00;
assign _c_characterGenerator[243] = 8'h18;
assign _c_characterGenerator[244] = 8'h18;
assign _c_characterGenerator[245] = 8'hdb;
assign _c_characterGenerator[246] = 8'h3c;
assign _c_characterGenerator[247] = 8'he7;
assign _c_characterGenerator[248] = 8'h3c;
assign _c_characterGenerator[249] = 8'hdb;
assign _c_characterGenerator[250] = 8'h18;
assign _c_characterGenerator[251] = 8'h18;
assign _c_characterGenerator[252] = 8'h00;
assign _c_characterGenerator[253] = 8'h00;
assign _c_characterGenerator[254] = 8'h00;
assign _c_characterGenerator[255] = 8'h00;
assign _c_characterGenerator[256] = 8'h00;
assign _c_characterGenerator[257] = 8'h80;
assign _c_characterGenerator[258] = 8'hc0;
assign _c_characterGenerator[259] = 8'he0;
assign _c_characterGenerator[260] = 8'hf0;
assign _c_characterGenerator[261] = 8'hf8;
assign _c_characterGenerator[262] = 8'hfe;
assign _c_characterGenerator[263] = 8'hf8;
assign _c_characterGenerator[264] = 8'hf0;
assign _c_characterGenerator[265] = 8'he0;
assign _c_characterGenerator[266] = 8'hc0;
assign _c_characterGenerator[267] = 8'h80;
assign _c_characterGenerator[268] = 8'h00;
assign _c_characterGenerator[269] = 8'h00;
assign _c_characterGenerator[270] = 8'h00;
assign _c_characterGenerator[271] = 8'h00;
assign _c_characterGenerator[272] = 8'h00;
assign _c_characterGenerator[273] = 8'h02;
assign _c_characterGenerator[274] = 8'h06;
assign _c_characterGenerator[275] = 8'h0e;
assign _c_characterGenerator[276] = 8'h1e;
assign _c_characterGenerator[277] = 8'h3e;
assign _c_characterGenerator[278] = 8'hfe;
assign _c_characterGenerator[279] = 8'h3e;
assign _c_characterGenerator[280] = 8'h1e;
assign _c_characterGenerator[281] = 8'h0e;
assign _c_characterGenerator[282] = 8'h06;
assign _c_characterGenerator[283] = 8'h02;
assign _c_characterGenerator[284] = 8'h00;
assign _c_characterGenerator[285] = 8'h00;
assign _c_characterGenerator[286] = 8'h00;
assign _c_characterGenerator[287] = 8'h00;
assign _c_characterGenerator[288] = 8'h00;
assign _c_characterGenerator[289] = 8'h00;
assign _c_characterGenerator[290] = 8'h18;
assign _c_characterGenerator[291] = 8'h3c;
assign _c_characterGenerator[292] = 8'h7e;
assign _c_characterGenerator[293] = 8'h18;
assign _c_characterGenerator[294] = 8'h18;
assign _c_characterGenerator[295] = 8'h18;
assign _c_characterGenerator[296] = 8'h7e;
assign _c_characterGenerator[297] = 8'h3c;
assign _c_characterGenerator[298] = 8'h18;
assign _c_characterGenerator[299] = 8'h00;
assign _c_characterGenerator[300] = 8'h00;
assign _c_characterGenerator[301] = 8'h00;
assign _c_characterGenerator[302] = 8'h00;
assign _c_characterGenerator[303] = 8'h00;
assign _c_characterGenerator[304] = 8'h00;
assign _c_characterGenerator[305] = 8'h00;
assign _c_characterGenerator[306] = 8'h66;
assign _c_characterGenerator[307] = 8'h66;
assign _c_characterGenerator[308] = 8'h66;
assign _c_characterGenerator[309] = 8'h66;
assign _c_characterGenerator[310] = 8'h66;
assign _c_characterGenerator[311] = 8'h66;
assign _c_characterGenerator[312] = 8'h66;
assign _c_characterGenerator[313] = 8'h00;
assign _c_characterGenerator[314] = 8'h66;
assign _c_characterGenerator[315] = 8'h66;
assign _c_characterGenerator[316] = 8'h00;
assign _c_characterGenerator[317] = 8'h00;
assign _c_characterGenerator[318] = 8'h00;
assign _c_characterGenerator[319] = 8'h00;
assign _c_characterGenerator[320] = 8'h00;
assign _c_characterGenerator[321] = 8'h00;
assign _c_characterGenerator[322] = 8'h7f;
assign _c_characterGenerator[323] = 8'hdb;
assign _c_characterGenerator[324] = 8'hdb;
assign _c_characterGenerator[325] = 8'hdb;
assign _c_characterGenerator[326] = 8'h7b;
assign _c_characterGenerator[327] = 8'h1b;
assign _c_characterGenerator[328] = 8'h1b;
assign _c_characterGenerator[329] = 8'h1b;
assign _c_characterGenerator[330] = 8'h1b;
assign _c_characterGenerator[331] = 8'h1b;
assign _c_characterGenerator[332] = 8'h00;
assign _c_characterGenerator[333] = 8'h00;
assign _c_characterGenerator[334] = 8'h00;
assign _c_characterGenerator[335] = 8'h00;
assign _c_characterGenerator[336] = 8'h00;
assign _c_characterGenerator[337] = 8'h7c;
assign _c_characterGenerator[338] = 8'hc6;
assign _c_characterGenerator[339] = 8'h60;
assign _c_characterGenerator[340] = 8'h38;
assign _c_characterGenerator[341] = 8'h6c;
assign _c_characterGenerator[342] = 8'hc6;
assign _c_characterGenerator[343] = 8'hc6;
assign _c_characterGenerator[344] = 8'h6c;
assign _c_characterGenerator[345] = 8'h38;
assign _c_characterGenerator[346] = 8'h0c;
assign _c_characterGenerator[347] = 8'hc6;
assign _c_characterGenerator[348] = 8'h7c;
assign _c_characterGenerator[349] = 8'h00;
assign _c_characterGenerator[350] = 8'h00;
assign _c_characterGenerator[351] = 8'h00;
assign _c_characterGenerator[352] = 8'h00;
assign _c_characterGenerator[353] = 8'h00;
assign _c_characterGenerator[354] = 8'h00;
assign _c_characterGenerator[355] = 8'h00;
assign _c_characterGenerator[356] = 8'h00;
assign _c_characterGenerator[357] = 8'h00;
assign _c_characterGenerator[358] = 8'h00;
assign _c_characterGenerator[359] = 8'h00;
assign _c_characterGenerator[360] = 8'hfe;
assign _c_characterGenerator[361] = 8'hfe;
assign _c_characterGenerator[362] = 8'hfe;
assign _c_characterGenerator[363] = 8'hfe;
assign _c_characterGenerator[364] = 8'h00;
assign _c_characterGenerator[365] = 8'h00;
assign _c_characterGenerator[366] = 8'h00;
assign _c_characterGenerator[367] = 8'h00;
assign _c_characterGenerator[368] = 8'h00;
assign _c_characterGenerator[369] = 8'h00;
assign _c_characterGenerator[370] = 8'h18;
assign _c_characterGenerator[371] = 8'h3c;
assign _c_characterGenerator[372] = 8'h7e;
assign _c_characterGenerator[373] = 8'h18;
assign _c_characterGenerator[374] = 8'h18;
assign _c_characterGenerator[375] = 8'h18;
assign _c_characterGenerator[376] = 8'h7e;
assign _c_characterGenerator[377] = 8'h3c;
assign _c_characterGenerator[378] = 8'h18;
assign _c_characterGenerator[379] = 8'h7e;
assign _c_characterGenerator[380] = 8'h00;
assign _c_characterGenerator[381] = 8'h00;
assign _c_characterGenerator[382] = 8'h00;
assign _c_characterGenerator[383] = 8'h00;
assign _c_characterGenerator[384] = 8'h00;
assign _c_characterGenerator[385] = 8'h00;
assign _c_characterGenerator[386] = 8'h18;
assign _c_characterGenerator[387] = 8'h3c;
assign _c_characterGenerator[388] = 8'h7e;
assign _c_characterGenerator[389] = 8'h18;
assign _c_characterGenerator[390] = 8'h18;
assign _c_characterGenerator[391] = 8'h18;
assign _c_characterGenerator[392] = 8'h18;
assign _c_characterGenerator[393] = 8'h18;
assign _c_characterGenerator[394] = 8'h18;
assign _c_characterGenerator[395] = 8'h18;
assign _c_characterGenerator[396] = 8'h00;
assign _c_characterGenerator[397] = 8'h00;
assign _c_characterGenerator[398] = 8'h00;
assign _c_characterGenerator[399] = 8'h00;
assign _c_characterGenerator[400] = 8'h00;
assign _c_characterGenerator[401] = 8'h00;
assign _c_characterGenerator[402] = 8'h18;
assign _c_characterGenerator[403] = 8'h18;
assign _c_characterGenerator[404] = 8'h18;
assign _c_characterGenerator[405] = 8'h18;
assign _c_characterGenerator[406] = 8'h18;
assign _c_characterGenerator[407] = 8'h18;
assign _c_characterGenerator[408] = 8'h18;
assign _c_characterGenerator[409] = 8'h7e;
assign _c_characterGenerator[410] = 8'h3c;
assign _c_characterGenerator[411] = 8'h18;
assign _c_characterGenerator[412] = 8'h00;
assign _c_characterGenerator[413] = 8'h00;
assign _c_characterGenerator[414] = 8'h00;
assign _c_characterGenerator[415] = 8'h00;
assign _c_characterGenerator[416] = 8'h00;
assign _c_characterGenerator[417] = 8'h00;
assign _c_characterGenerator[418] = 8'h00;
assign _c_characterGenerator[419] = 8'h00;
assign _c_characterGenerator[420] = 8'h00;
assign _c_characterGenerator[421] = 8'h18;
assign _c_characterGenerator[422] = 8'h0c;
assign _c_characterGenerator[423] = 8'hfe;
assign _c_characterGenerator[424] = 8'h0c;
assign _c_characterGenerator[425] = 8'h18;
assign _c_characterGenerator[426] = 8'h00;
assign _c_characterGenerator[427] = 8'h00;
assign _c_characterGenerator[428] = 8'h00;
assign _c_characterGenerator[429] = 8'h00;
assign _c_characterGenerator[430] = 8'h00;
assign _c_characterGenerator[431] = 8'h00;
assign _c_characterGenerator[432] = 8'h00;
assign _c_characterGenerator[433] = 8'h00;
assign _c_characterGenerator[434] = 8'h00;
assign _c_characterGenerator[435] = 8'h00;
assign _c_characterGenerator[436] = 8'h00;
assign _c_characterGenerator[437] = 8'h30;
assign _c_characterGenerator[438] = 8'h60;
assign _c_characterGenerator[439] = 8'hfe;
assign _c_characterGenerator[440] = 8'h60;
assign _c_characterGenerator[441] = 8'h30;
assign _c_characterGenerator[442] = 8'h00;
assign _c_characterGenerator[443] = 8'h00;
assign _c_characterGenerator[444] = 8'h00;
assign _c_characterGenerator[445] = 8'h00;
assign _c_characterGenerator[446] = 8'h00;
assign _c_characterGenerator[447] = 8'h00;
assign _c_characterGenerator[448] = 8'h00;
assign _c_characterGenerator[449] = 8'h00;
assign _c_characterGenerator[450] = 8'h00;
assign _c_characterGenerator[451] = 8'h00;
assign _c_characterGenerator[452] = 8'h00;
assign _c_characterGenerator[453] = 8'h00;
assign _c_characterGenerator[454] = 8'hc0;
assign _c_characterGenerator[455] = 8'hc0;
assign _c_characterGenerator[456] = 8'hc0;
assign _c_characterGenerator[457] = 8'hfe;
assign _c_characterGenerator[458] = 8'h00;
assign _c_characterGenerator[459] = 8'h00;
assign _c_characterGenerator[460] = 8'h00;
assign _c_characterGenerator[461] = 8'h00;
assign _c_characterGenerator[462] = 8'h00;
assign _c_characterGenerator[463] = 8'h00;
assign _c_characterGenerator[464] = 8'h00;
assign _c_characterGenerator[465] = 8'h00;
assign _c_characterGenerator[466] = 8'h00;
assign _c_characterGenerator[467] = 8'h00;
assign _c_characterGenerator[468] = 8'h00;
assign _c_characterGenerator[469] = 8'h28;
assign _c_characterGenerator[470] = 8'h6c;
assign _c_characterGenerator[471] = 8'hfe;
assign _c_characterGenerator[472] = 8'h6c;
assign _c_characterGenerator[473] = 8'h28;
assign _c_characterGenerator[474] = 8'h00;
assign _c_characterGenerator[475] = 8'h00;
assign _c_characterGenerator[476] = 8'h00;
assign _c_characterGenerator[477] = 8'h00;
assign _c_characterGenerator[478] = 8'h00;
assign _c_characterGenerator[479] = 8'h00;
assign _c_characterGenerator[480] = 8'h00;
assign _c_characterGenerator[481] = 8'h00;
assign _c_characterGenerator[482] = 8'h00;
assign _c_characterGenerator[483] = 8'h00;
assign _c_characterGenerator[484] = 8'h10;
assign _c_characterGenerator[485] = 8'h38;
assign _c_characterGenerator[486] = 8'h38;
assign _c_characterGenerator[487] = 8'h7c;
assign _c_characterGenerator[488] = 8'h7c;
assign _c_characterGenerator[489] = 8'hfe;
assign _c_characterGenerator[490] = 8'hfe;
assign _c_characterGenerator[491] = 8'h00;
assign _c_characterGenerator[492] = 8'h00;
assign _c_characterGenerator[493] = 8'h00;
assign _c_characterGenerator[494] = 8'h00;
assign _c_characterGenerator[495] = 8'h00;
assign _c_characterGenerator[496] = 8'h00;
assign _c_characterGenerator[497] = 8'h00;
assign _c_characterGenerator[498] = 8'h00;
assign _c_characterGenerator[499] = 8'h00;
assign _c_characterGenerator[500] = 8'hfe;
assign _c_characterGenerator[501] = 8'hfe;
assign _c_characterGenerator[502] = 8'h7c;
assign _c_characterGenerator[503] = 8'h7c;
assign _c_characterGenerator[504] = 8'h38;
assign _c_characterGenerator[505] = 8'h38;
assign _c_characterGenerator[506] = 8'h10;
assign _c_characterGenerator[507] = 8'h00;
assign _c_characterGenerator[508] = 8'h00;
assign _c_characterGenerator[509] = 8'h00;
assign _c_characterGenerator[510] = 8'h00;
assign _c_characterGenerator[511] = 8'h00;
assign _c_characterGenerator[512] = 8'h00;
assign _c_characterGenerator[513] = 8'h00;
assign _c_characterGenerator[514] = 8'h00;
assign _c_characterGenerator[515] = 8'h00;
assign _c_characterGenerator[516] = 8'h00;
assign _c_characterGenerator[517] = 8'h00;
assign _c_characterGenerator[518] = 8'h00;
assign _c_characterGenerator[519] = 8'h00;
assign _c_characterGenerator[520] = 8'h00;
assign _c_characterGenerator[521] = 8'h00;
assign _c_characterGenerator[522] = 8'h00;
assign _c_characterGenerator[523] = 8'h00;
assign _c_characterGenerator[524] = 8'h00;
assign _c_characterGenerator[525] = 8'h00;
assign _c_characterGenerator[526] = 8'h00;
assign _c_characterGenerator[527] = 8'h00;
assign _c_characterGenerator[528] = 8'h00;
assign _c_characterGenerator[529] = 8'h00;
assign _c_characterGenerator[530] = 8'h18;
assign _c_characterGenerator[531] = 8'h3c;
assign _c_characterGenerator[532] = 8'h3c;
assign _c_characterGenerator[533] = 8'h3c;
assign _c_characterGenerator[534] = 8'h18;
assign _c_characterGenerator[535] = 8'h18;
assign _c_characterGenerator[536] = 8'h18;
assign _c_characterGenerator[537] = 8'h00;
assign _c_characterGenerator[538] = 8'h18;
assign _c_characterGenerator[539] = 8'h18;
assign _c_characterGenerator[540] = 8'h00;
assign _c_characterGenerator[541] = 8'h00;
assign _c_characterGenerator[542] = 8'h00;
assign _c_characterGenerator[543] = 8'h00;
assign _c_characterGenerator[544] = 8'h00;
assign _c_characterGenerator[545] = 8'h66;
assign _c_characterGenerator[546] = 8'h66;
assign _c_characterGenerator[547] = 8'h66;
assign _c_characterGenerator[548] = 8'h24;
assign _c_characterGenerator[549] = 8'h00;
assign _c_characterGenerator[550] = 8'h00;
assign _c_characterGenerator[551] = 8'h00;
assign _c_characterGenerator[552] = 8'h00;
assign _c_characterGenerator[553] = 8'h00;
assign _c_characterGenerator[554] = 8'h00;
assign _c_characterGenerator[555] = 8'h00;
assign _c_characterGenerator[556] = 8'h00;
assign _c_characterGenerator[557] = 8'h00;
assign _c_characterGenerator[558] = 8'h00;
assign _c_characterGenerator[559] = 8'h00;
assign _c_characterGenerator[560] = 8'h00;
assign _c_characterGenerator[561] = 8'h00;
assign _c_characterGenerator[562] = 8'h00;
assign _c_characterGenerator[563] = 8'h6c;
assign _c_characterGenerator[564] = 8'h6c;
assign _c_characterGenerator[565] = 8'hfe;
assign _c_characterGenerator[566] = 8'h6c;
assign _c_characterGenerator[567] = 8'h6c;
assign _c_characterGenerator[568] = 8'h6c;
assign _c_characterGenerator[569] = 8'hfe;
assign _c_characterGenerator[570] = 8'h6c;
assign _c_characterGenerator[571] = 8'h6c;
assign _c_characterGenerator[572] = 8'h00;
assign _c_characterGenerator[573] = 8'h00;
assign _c_characterGenerator[574] = 8'h00;
assign _c_characterGenerator[575] = 8'h00;
assign _c_characterGenerator[576] = 8'h18;
assign _c_characterGenerator[577] = 8'h18;
assign _c_characterGenerator[578] = 8'h7c;
assign _c_characterGenerator[579] = 8'hc6;
assign _c_characterGenerator[580] = 8'hc2;
assign _c_characterGenerator[581] = 8'hc0;
assign _c_characterGenerator[582] = 8'h7c;
assign _c_characterGenerator[583] = 8'h06;
assign _c_characterGenerator[584] = 8'h06;
assign _c_characterGenerator[585] = 8'h86;
assign _c_characterGenerator[586] = 8'hc6;
assign _c_characterGenerator[587] = 8'h7c;
assign _c_characterGenerator[588] = 8'h18;
assign _c_characterGenerator[589] = 8'h18;
assign _c_characterGenerator[590] = 8'h00;
assign _c_characterGenerator[591] = 8'h00;
assign _c_characterGenerator[592] = 8'h00;
assign _c_characterGenerator[593] = 8'h00;
assign _c_characterGenerator[594] = 8'h00;
assign _c_characterGenerator[595] = 8'h00;
assign _c_characterGenerator[596] = 8'hc2;
assign _c_characterGenerator[597] = 8'hc6;
assign _c_characterGenerator[598] = 8'h0c;
assign _c_characterGenerator[599] = 8'h18;
assign _c_characterGenerator[600] = 8'h30;
assign _c_characterGenerator[601] = 8'h60;
assign _c_characterGenerator[602] = 8'hc6;
assign _c_characterGenerator[603] = 8'h86;
assign _c_characterGenerator[604] = 8'h00;
assign _c_characterGenerator[605] = 8'h00;
assign _c_characterGenerator[606] = 8'h00;
assign _c_characterGenerator[607] = 8'h00;
assign _c_characterGenerator[608] = 8'h00;
assign _c_characterGenerator[609] = 8'h00;
assign _c_characterGenerator[610] = 8'h38;
assign _c_characterGenerator[611] = 8'h6c;
assign _c_characterGenerator[612] = 8'h6c;
assign _c_characterGenerator[613] = 8'h38;
assign _c_characterGenerator[614] = 8'h76;
assign _c_characterGenerator[615] = 8'hdc;
assign _c_characterGenerator[616] = 8'hcc;
assign _c_characterGenerator[617] = 8'hcc;
assign _c_characterGenerator[618] = 8'hcc;
assign _c_characterGenerator[619] = 8'h76;
assign _c_characterGenerator[620] = 8'h00;
assign _c_characterGenerator[621] = 8'h00;
assign _c_characterGenerator[622] = 8'h00;
assign _c_characterGenerator[623] = 8'h00;
assign _c_characterGenerator[624] = 8'h00;
assign _c_characterGenerator[625] = 8'h30;
assign _c_characterGenerator[626] = 8'h30;
assign _c_characterGenerator[627] = 8'h30;
assign _c_characterGenerator[628] = 8'h60;
assign _c_characterGenerator[629] = 8'h00;
assign _c_characterGenerator[630] = 8'h00;
assign _c_characterGenerator[631] = 8'h00;
assign _c_characterGenerator[632] = 8'h00;
assign _c_characterGenerator[633] = 8'h00;
assign _c_characterGenerator[634] = 8'h00;
assign _c_characterGenerator[635] = 8'h00;
assign _c_characterGenerator[636] = 8'h00;
assign _c_characterGenerator[637] = 8'h00;
assign _c_characterGenerator[638] = 8'h00;
assign _c_characterGenerator[639] = 8'h00;
assign _c_characterGenerator[640] = 8'h00;
assign _c_characterGenerator[641] = 8'h00;
assign _c_characterGenerator[642] = 8'h0c;
assign _c_characterGenerator[643] = 8'h18;
assign _c_characterGenerator[644] = 8'h30;
assign _c_characterGenerator[645] = 8'h30;
assign _c_characterGenerator[646] = 8'h30;
assign _c_characterGenerator[647] = 8'h30;
assign _c_characterGenerator[648] = 8'h30;
assign _c_characterGenerator[649] = 8'h30;
assign _c_characterGenerator[650] = 8'h18;
assign _c_characterGenerator[651] = 8'h0c;
assign _c_characterGenerator[652] = 8'h00;
assign _c_characterGenerator[653] = 8'h00;
assign _c_characterGenerator[654] = 8'h00;
assign _c_characterGenerator[655] = 8'h00;
assign _c_characterGenerator[656] = 8'h00;
assign _c_characterGenerator[657] = 8'h00;
assign _c_characterGenerator[658] = 8'h30;
assign _c_characterGenerator[659] = 8'h18;
assign _c_characterGenerator[660] = 8'h0c;
assign _c_characterGenerator[661] = 8'h0c;
assign _c_characterGenerator[662] = 8'h0c;
assign _c_characterGenerator[663] = 8'h0c;
assign _c_characterGenerator[664] = 8'h0c;
assign _c_characterGenerator[665] = 8'h0c;
assign _c_characterGenerator[666] = 8'h18;
assign _c_characterGenerator[667] = 8'h30;
assign _c_characterGenerator[668] = 8'h00;
assign _c_characterGenerator[669] = 8'h00;
assign _c_characterGenerator[670] = 8'h00;
assign _c_characterGenerator[671] = 8'h00;
assign _c_characterGenerator[672] = 8'h00;
assign _c_characterGenerator[673] = 8'h00;
assign _c_characterGenerator[674] = 8'h00;
assign _c_characterGenerator[675] = 8'h00;
assign _c_characterGenerator[676] = 8'h00;
assign _c_characterGenerator[677] = 8'h66;
assign _c_characterGenerator[678] = 8'h3c;
assign _c_characterGenerator[679] = 8'hff;
assign _c_characterGenerator[680] = 8'h3c;
assign _c_characterGenerator[681] = 8'h66;
assign _c_characterGenerator[682] = 8'h00;
assign _c_characterGenerator[683] = 8'h00;
assign _c_characterGenerator[684] = 8'h00;
assign _c_characterGenerator[685] = 8'h00;
assign _c_characterGenerator[686] = 8'h00;
assign _c_characterGenerator[687] = 8'h00;
assign _c_characterGenerator[688] = 8'h00;
assign _c_characterGenerator[689] = 8'h00;
assign _c_characterGenerator[690] = 8'h00;
assign _c_characterGenerator[691] = 8'h00;
assign _c_characterGenerator[692] = 8'h00;
assign _c_characterGenerator[693] = 8'h18;
assign _c_characterGenerator[694] = 8'h18;
assign _c_characterGenerator[695] = 8'h7e;
assign _c_characterGenerator[696] = 8'h18;
assign _c_characterGenerator[697] = 8'h18;
assign _c_characterGenerator[698] = 8'h00;
assign _c_characterGenerator[699] = 8'h00;
assign _c_characterGenerator[700] = 8'h00;
assign _c_characterGenerator[701] = 8'h00;
assign _c_characterGenerator[702] = 8'h00;
assign _c_characterGenerator[703] = 8'h00;
assign _c_characterGenerator[704] = 8'h00;
assign _c_characterGenerator[705] = 8'h00;
assign _c_characterGenerator[706] = 8'h00;
assign _c_characterGenerator[707] = 8'h00;
assign _c_characterGenerator[708] = 8'h00;
assign _c_characterGenerator[709] = 8'h00;
assign _c_characterGenerator[710] = 8'h00;
assign _c_characterGenerator[711] = 8'h00;
assign _c_characterGenerator[712] = 8'h00;
assign _c_characterGenerator[713] = 8'h18;
assign _c_characterGenerator[714] = 8'h18;
assign _c_characterGenerator[715] = 8'h18;
assign _c_characterGenerator[716] = 8'h30;
assign _c_characterGenerator[717] = 8'h00;
assign _c_characterGenerator[718] = 8'h00;
assign _c_characterGenerator[719] = 8'h00;
assign _c_characterGenerator[720] = 8'h00;
assign _c_characterGenerator[721] = 8'h00;
assign _c_characterGenerator[722] = 8'h00;
assign _c_characterGenerator[723] = 8'h00;
assign _c_characterGenerator[724] = 8'h00;
assign _c_characterGenerator[725] = 8'h00;
assign _c_characterGenerator[726] = 8'h00;
assign _c_characterGenerator[727] = 8'hfe;
assign _c_characterGenerator[728] = 8'h00;
assign _c_characterGenerator[729] = 8'h00;
assign _c_characterGenerator[730] = 8'h00;
assign _c_characterGenerator[731] = 8'h00;
assign _c_characterGenerator[732] = 8'h00;
assign _c_characterGenerator[733] = 8'h00;
assign _c_characterGenerator[734] = 8'h00;
assign _c_characterGenerator[735] = 8'h00;
assign _c_characterGenerator[736] = 8'h00;
assign _c_characterGenerator[737] = 8'h00;
assign _c_characterGenerator[738] = 8'h00;
assign _c_characterGenerator[739] = 8'h00;
assign _c_characterGenerator[740] = 8'h00;
assign _c_characterGenerator[741] = 8'h00;
assign _c_characterGenerator[742] = 8'h00;
assign _c_characterGenerator[743] = 8'h00;
assign _c_characterGenerator[744] = 8'h00;
assign _c_characterGenerator[745] = 8'h00;
assign _c_characterGenerator[746] = 8'h18;
assign _c_characterGenerator[747] = 8'h18;
assign _c_characterGenerator[748] = 8'h00;
assign _c_characterGenerator[749] = 8'h00;
assign _c_characterGenerator[750] = 8'h00;
assign _c_characterGenerator[751] = 8'h00;
assign _c_characterGenerator[752] = 8'h00;
assign _c_characterGenerator[753] = 8'h00;
assign _c_characterGenerator[754] = 8'h00;
assign _c_characterGenerator[755] = 8'h00;
assign _c_characterGenerator[756] = 8'h02;
assign _c_characterGenerator[757] = 8'h06;
assign _c_characterGenerator[758] = 8'h0c;
assign _c_characterGenerator[759] = 8'h18;
assign _c_characterGenerator[760] = 8'h30;
assign _c_characterGenerator[761] = 8'h60;
assign _c_characterGenerator[762] = 8'hc0;
assign _c_characterGenerator[763] = 8'h80;
assign _c_characterGenerator[764] = 8'h00;
assign _c_characterGenerator[765] = 8'h00;
assign _c_characterGenerator[766] = 8'h00;
assign _c_characterGenerator[767] = 8'h00;
assign _c_characterGenerator[768] = 8'h00;
assign _c_characterGenerator[769] = 8'h00;
assign _c_characterGenerator[770] = 8'h38;
assign _c_characterGenerator[771] = 8'h6c;
assign _c_characterGenerator[772] = 8'hc6;
assign _c_characterGenerator[773] = 8'hc6;
assign _c_characterGenerator[774] = 8'hd6;
assign _c_characterGenerator[775] = 8'hd6;
assign _c_characterGenerator[776] = 8'hc6;
assign _c_characterGenerator[777] = 8'hc6;
assign _c_characterGenerator[778] = 8'h6c;
assign _c_characterGenerator[779] = 8'h38;
assign _c_characterGenerator[780] = 8'h00;
assign _c_characterGenerator[781] = 8'h00;
assign _c_characterGenerator[782] = 8'h00;
assign _c_characterGenerator[783] = 8'h00;
assign _c_characterGenerator[784] = 8'h00;
assign _c_characterGenerator[785] = 8'h00;
assign _c_characterGenerator[786] = 8'h18;
assign _c_characterGenerator[787] = 8'h38;
assign _c_characterGenerator[788] = 8'h78;
assign _c_characterGenerator[789] = 8'h18;
assign _c_characterGenerator[790] = 8'h18;
assign _c_characterGenerator[791] = 8'h18;
assign _c_characterGenerator[792] = 8'h18;
assign _c_characterGenerator[793] = 8'h18;
assign _c_characterGenerator[794] = 8'h18;
assign _c_characterGenerator[795] = 8'h7e;
assign _c_characterGenerator[796] = 8'h00;
assign _c_characterGenerator[797] = 8'h00;
assign _c_characterGenerator[798] = 8'h00;
assign _c_characterGenerator[799] = 8'h00;
assign _c_characterGenerator[800] = 8'h00;
assign _c_characterGenerator[801] = 8'h00;
assign _c_characterGenerator[802] = 8'h7c;
assign _c_characterGenerator[803] = 8'hc6;
assign _c_characterGenerator[804] = 8'h06;
assign _c_characterGenerator[805] = 8'h0c;
assign _c_characterGenerator[806] = 8'h18;
assign _c_characterGenerator[807] = 8'h30;
assign _c_characterGenerator[808] = 8'h60;
assign _c_characterGenerator[809] = 8'hc0;
assign _c_characterGenerator[810] = 8'hc6;
assign _c_characterGenerator[811] = 8'hfe;
assign _c_characterGenerator[812] = 8'h00;
assign _c_characterGenerator[813] = 8'h00;
assign _c_characterGenerator[814] = 8'h00;
assign _c_characterGenerator[815] = 8'h00;
assign _c_characterGenerator[816] = 8'h00;
assign _c_characterGenerator[817] = 8'h00;
assign _c_characterGenerator[818] = 8'h7c;
assign _c_characterGenerator[819] = 8'hc6;
assign _c_characterGenerator[820] = 8'h06;
assign _c_characterGenerator[821] = 8'h06;
assign _c_characterGenerator[822] = 8'h3c;
assign _c_characterGenerator[823] = 8'h06;
assign _c_characterGenerator[824] = 8'h06;
assign _c_characterGenerator[825] = 8'h06;
assign _c_characterGenerator[826] = 8'hc6;
assign _c_characterGenerator[827] = 8'h7c;
assign _c_characterGenerator[828] = 8'h00;
assign _c_characterGenerator[829] = 8'h00;
assign _c_characterGenerator[830] = 8'h00;
assign _c_characterGenerator[831] = 8'h00;
assign _c_characterGenerator[832] = 8'h00;
assign _c_characterGenerator[833] = 8'h00;
assign _c_characterGenerator[834] = 8'h0c;
assign _c_characterGenerator[835] = 8'h1c;
assign _c_characterGenerator[836] = 8'h3c;
assign _c_characterGenerator[837] = 8'h6c;
assign _c_characterGenerator[838] = 8'hcc;
assign _c_characterGenerator[839] = 8'hfe;
assign _c_characterGenerator[840] = 8'h0c;
assign _c_characterGenerator[841] = 8'h0c;
assign _c_characterGenerator[842] = 8'h0c;
assign _c_characterGenerator[843] = 8'h1e;
assign _c_characterGenerator[844] = 8'h00;
assign _c_characterGenerator[845] = 8'h00;
assign _c_characterGenerator[846] = 8'h00;
assign _c_characterGenerator[847] = 8'h00;
assign _c_characterGenerator[848] = 8'h00;
assign _c_characterGenerator[849] = 8'h00;
assign _c_characterGenerator[850] = 8'hfe;
assign _c_characterGenerator[851] = 8'hc0;
assign _c_characterGenerator[852] = 8'hc0;
assign _c_characterGenerator[853] = 8'hc0;
assign _c_characterGenerator[854] = 8'hfc;
assign _c_characterGenerator[855] = 8'h06;
assign _c_characterGenerator[856] = 8'h06;
assign _c_characterGenerator[857] = 8'h06;
assign _c_characterGenerator[858] = 8'hc6;
assign _c_characterGenerator[859] = 8'h7c;
assign _c_characterGenerator[860] = 8'h00;
assign _c_characterGenerator[861] = 8'h00;
assign _c_characterGenerator[862] = 8'h00;
assign _c_characterGenerator[863] = 8'h00;
assign _c_characterGenerator[864] = 8'h00;
assign _c_characterGenerator[865] = 8'h00;
assign _c_characterGenerator[866] = 8'h38;
assign _c_characterGenerator[867] = 8'h60;
assign _c_characterGenerator[868] = 8'hc0;
assign _c_characterGenerator[869] = 8'hc0;
assign _c_characterGenerator[870] = 8'hfc;
assign _c_characterGenerator[871] = 8'hc6;
assign _c_characterGenerator[872] = 8'hc6;
assign _c_characterGenerator[873] = 8'hc6;
assign _c_characterGenerator[874] = 8'hc6;
assign _c_characterGenerator[875] = 8'h7c;
assign _c_characterGenerator[876] = 8'h00;
assign _c_characterGenerator[877] = 8'h00;
assign _c_characterGenerator[878] = 8'h00;
assign _c_characterGenerator[879] = 8'h00;
assign _c_characterGenerator[880] = 8'h00;
assign _c_characterGenerator[881] = 8'h00;
assign _c_characterGenerator[882] = 8'hfe;
assign _c_characterGenerator[883] = 8'hc6;
assign _c_characterGenerator[884] = 8'h06;
assign _c_characterGenerator[885] = 8'h06;
assign _c_characterGenerator[886] = 8'h0c;
assign _c_characterGenerator[887] = 8'h18;
assign _c_characterGenerator[888] = 8'h30;
assign _c_characterGenerator[889] = 8'h30;
assign _c_characterGenerator[890] = 8'h30;
assign _c_characterGenerator[891] = 8'h30;
assign _c_characterGenerator[892] = 8'h00;
assign _c_characterGenerator[893] = 8'h00;
assign _c_characterGenerator[894] = 8'h00;
assign _c_characterGenerator[895] = 8'h00;
assign _c_characterGenerator[896] = 8'h00;
assign _c_characterGenerator[897] = 8'h00;
assign _c_characterGenerator[898] = 8'h7c;
assign _c_characterGenerator[899] = 8'hc6;
assign _c_characterGenerator[900] = 8'hc6;
assign _c_characterGenerator[901] = 8'hc6;
assign _c_characterGenerator[902] = 8'h7c;
assign _c_characterGenerator[903] = 8'hc6;
assign _c_characterGenerator[904] = 8'hc6;
assign _c_characterGenerator[905] = 8'hc6;
assign _c_characterGenerator[906] = 8'hc6;
assign _c_characterGenerator[907] = 8'h7c;
assign _c_characterGenerator[908] = 8'h00;
assign _c_characterGenerator[909] = 8'h00;
assign _c_characterGenerator[910] = 8'h00;
assign _c_characterGenerator[911] = 8'h00;
assign _c_characterGenerator[912] = 8'h00;
assign _c_characterGenerator[913] = 8'h00;
assign _c_characterGenerator[914] = 8'h7c;
assign _c_characterGenerator[915] = 8'hc6;
assign _c_characterGenerator[916] = 8'hc6;
assign _c_characterGenerator[917] = 8'hc6;
assign _c_characterGenerator[918] = 8'h7e;
assign _c_characterGenerator[919] = 8'h06;
assign _c_characterGenerator[920] = 8'h06;
assign _c_characterGenerator[921] = 8'h06;
assign _c_characterGenerator[922] = 8'h0c;
assign _c_characterGenerator[923] = 8'h78;
assign _c_characterGenerator[924] = 8'h00;
assign _c_characterGenerator[925] = 8'h00;
assign _c_characterGenerator[926] = 8'h00;
assign _c_characterGenerator[927] = 8'h00;
assign _c_characterGenerator[928] = 8'h00;
assign _c_characterGenerator[929] = 8'h00;
assign _c_characterGenerator[930] = 8'h00;
assign _c_characterGenerator[931] = 8'h00;
assign _c_characterGenerator[932] = 8'h18;
assign _c_characterGenerator[933] = 8'h18;
assign _c_characterGenerator[934] = 8'h00;
assign _c_characterGenerator[935] = 8'h00;
assign _c_characterGenerator[936] = 8'h00;
assign _c_characterGenerator[937] = 8'h18;
assign _c_characterGenerator[938] = 8'h18;
assign _c_characterGenerator[939] = 8'h00;
assign _c_characterGenerator[940] = 8'h00;
assign _c_characterGenerator[941] = 8'h00;
assign _c_characterGenerator[942] = 8'h00;
assign _c_characterGenerator[943] = 8'h00;
assign _c_characterGenerator[944] = 8'h00;
assign _c_characterGenerator[945] = 8'h00;
assign _c_characterGenerator[946] = 8'h00;
assign _c_characterGenerator[947] = 8'h00;
assign _c_characterGenerator[948] = 8'h18;
assign _c_characterGenerator[949] = 8'h18;
assign _c_characterGenerator[950] = 8'h00;
assign _c_characterGenerator[951] = 8'h00;
assign _c_characterGenerator[952] = 8'h00;
assign _c_characterGenerator[953] = 8'h18;
assign _c_characterGenerator[954] = 8'h18;
assign _c_characterGenerator[955] = 8'h30;
assign _c_characterGenerator[956] = 8'h00;
assign _c_characterGenerator[957] = 8'h00;
assign _c_characterGenerator[958] = 8'h00;
assign _c_characterGenerator[959] = 8'h00;
assign _c_characterGenerator[960] = 8'h00;
assign _c_characterGenerator[961] = 8'h00;
assign _c_characterGenerator[962] = 8'h00;
assign _c_characterGenerator[963] = 8'h06;
assign _c_characterGenerator[964] = 8'h0c;
assign _c_characterGenerator[965] = 8'h18;
assign _c_characterGenerator[966] = 8'h30;
assign _c_characterGenerator[967] = 8'h60;
assign _c_characterGenerator[968] = 8'h30;
assign _c_characterGenerator[969] = 8'h18;
assign _c_characterGenerator[970] = 8'h0c;
assign _c_characterGenerator[971] = 8'h06;
assign _c_characterGenerator[972] = 8'h00;
assign _c_characterGenerator[973] = 8'h00;
assign _c_characterGenerator[974] = 8'h00;
assign _c_characterGenerator[975] = 8'h00;
assign _c_characterGenerator[976] = 8'h00;
assign _c_characterGenerator[977] = 8'h00;
assign _c_characterGenerator[978] = 8'h00;
assign _c_characterGenerator[979] = 8'h00;
assign _c_characterGenerator[980] = 8'h00;
assign _c_characterGenerator[981] = 8'h7e;
assign _c_characterGenerator[982] = 8'h00;
assign _c_characterGenerator[983] = 8'h00;
assign _c_characterGenerator[984] = 8'h7e;
assign _c_characterGenerator[985] = 8'h00;
assign _c_characterGenerator[986] = 8'h00;
assign _c_characterGenerator[987] = 8'h00;
assign _c_characterGenerator[988] = 8'h00;
assign _c_characterGenerator[989] = 8'h00;
assign _c_characterGenerator[990] = 8'h00;
assign _c_characterGenerator[991] = 8'h00;
assign _c_characterGenerator[992] = 8'h00;
assign _c_characterGenerator[993] = 8'h00;
assign _c_characterGenerator[994] = 8'h00;
assign _c_characterGenerator[995] = 8'h60;
assign _c_characterGenerator[996] = 8'h30;
assign _c_characterGenerator[997] = 8'h18;
assign _c_characterGenerator[998] = 8'h0c;
assign _c_characterGenerator[999] = 8'h06;
assign _c_characterGenerator[1000] = 8'h0c;
assign _c_characterGenerator[1001] = 8'h18;
assign _c_characterGenerator[1002] = 8'h30;
assign _c_characterGenerator[1003] = 8'h60;
assign _c_characterGenerator[1004] = 8'h00;
assign _c_characterGenerator[1005] = 8'h00;
assign _c_characterGenerator[1006] = 8'h00;
assign _c_characterGenerator[1007] = 8'h00;
assign _c_characterGenerator[1008] = 8'h00;
assign _c_characterGenerator[1009] = 8'h00;
assign _c_characterGenerator[1010] = 8'h7c;
assign _c_characterGenerator[1011] = 8'hc6;
assign _c_characterGenerator[1012] = 8'hc6;
assign _c_characterGenerator[1013] = 8'h0c;
assign _c_characterGenerator[1014] = 8'h18;
assign _c_characterGenerator[1015] = 8'h18;
assign _c_characterGenerator[1016] = 8'h18;
assign _c_characterGenerator[1017] = 8'h00;
assign _c_characterGenerator[1018] = 8'h18;
assign _c_characterGenerator[1019] = 8'h18;
assign _c_characterGenerator[1020] = 8'h00;
assign _c_characterGenerator[1021] = 8'h00;
assign _c_characterGenerator[1022] = 8'h00;
assign _c_characterGenerator[1023] = 8'h00;
assign _c_characterGenerator[1024] = 8'h00;
assign _c_characterGenerator[1025] = 8'h00;
assign _c_characterGenerator[1026] = 8'h00;
assign _c_characterGenerator[1027] = 8'h7c;
assign _c_characterGenerator[1028] = 8'hc6;
assign _c_characterGenerator[1029] = 8'hc6;
assign _c_characterGenerator[1030] = 8'hde;
assign _c_characterGenerator[1031] = 8'hde;
assign _c_characterGenerator[1032] = 8'hde;
assign _c_characterGenerator[1033] = 8'hdc;
assign _c_characterGenerator[1034] = 8'hc0;
assign _c_characterGenerator[1035] = 8'h7c;
assign _c_characterGenerator[1036] = 8'h00;
assign _c_characterGenerator[1037] = 8'h00;
assign _c_characterGenerator[1038] = 8'h00;
assign _c_characterGenerator[1039] = 8'h00;
assign _c_characterGenerator[1040] = 8'h00;
assign _c_characterGenerator[1041] = 8'h00;
assign _c_characterGenerator[1042] = 8'h10;
assign _c_characterGenerator[1043] = 8'h38;
assign _c_characterGenerator[1044] = 8'h6c;
assign _c_characterGenerator[1045] = 8'hc6;
assign _c_characterGenerator[1046] = 8'hc6;
assign _c_characterGenerator[1047] = 8'hfe;
assign _c_characterGenerator[1048] = 8'hc6;
assign _c_characterGenerator[1049] = 8'hc6;
assign _c_characterGenerator[1050] = 8'hc6;
assign _c_characterGenerator[1051] = 8'hc6;
assign _c_characterGenerator[1052] = 8'h00;
assign _c_characterGenerator[1053] = 8'h00;
assign _c_characterGenerator[1054] = 8'h00;
assign _c_characterGenerator[1055] = 8'h00;
assign _c_characterGenerator[1056] = 8'h00;
assign _c_characterGenerator[1057] = 8'h00;
assign _c_characterGenerator[1058] = 8'hfc;
assign _c_characterGenerator[1059] = 8'h66;
assign _c_characterGenerator[1060] = 8'h66;
assign _c_characterGenerator[1061] = 8'h66;
assign _c_characterGenerator[1062] = 8'h7c;
assign _c_characterGenerator[1063] = 8'h66;
assign _c_characterGenerator[1064] = 8'h66;
assign _c_characterGenerator[1065] = 8'h66;
assign _c_characterGenerator[1066] = 8'h66;
assign _c_characterGenerator[1067] = 8'hfc;
assign _c_characterGenerator[1068] = 8'h00;
assign _c_characterGenerator[1069] = 8'h00;
assign _c_characterGenerator[1070] = 8'h00;
assign _c_characterGenerator[1071] = 8'h00;
assign _c_characterGenerator[1072] = 8'h00;
assign _c_characterGenerator[1073] = 8'h00;
assign _c_characterGenerator[1074] = 8'h3c;
assign _c_characterGenerator[1075] = 8'h66;
assign _c_characterGenerator[1076] = 8'hc2;
assign _c_characterGenerator[1077] = 8'hc0;
assign _c_characterGenerator[1078] = 8'hc0;
assign _c_characterGenerator[1079] = 8'hc0;
assign _c_characterGenerator[1080] = 8'hc0;
assign _c_characterGenerator[1081] = 8'hc2;
assign _c_characterGenerator[1082] = 8'h66;
assign _c_characterGenerator[1083] = 8'h3c;
assign _c_characterGenerator[1084] = 8'h00;
assign _c_characterGenerator[1085] = 8'h00;
assign _c_characterGenerator[1086] = 8'h00;
assign _c_characterGenerator[1087] = 8'h00;
assign _c_characterGenerator[1088] = 8'h00;
assign _c_characterGenerator[1089] = 8'h00;
assign _c_characterGenerator[1090] = 8'hf8;
assign _c_characterGenerator[1091] = 8'h6c;
assign _c_characterGenerator[1092] = 8'h66;
assign _c_characterGenerator[1093] = 8'h66;
assign _c_characterGenerator[1094] = 8'h66;
assign _c_characterGenerator[1095] = 8'h66;
assign _c_characterGenerator[1096] = 8'h66;
assign _c_characterGenerator[1097] = 8'h66;
assign _c_characterGenerator[1098] = 8'h6c;
assign _c_characterGenerator[1099] = 8'hf8;
assign _c_characterGenerator[1100] = 8'h00;
assign _c_characterGenerator[1101] = 8'h00;
assign _c_characterGenerator[1102] = 8'h00;
assign _c_characterGenerator[1103] = 8'h00;
assign _c_characterGenerator[1104] = 8'h00;
assign _c_characterGenerator[1105] = 8'h00;
assign _c_characterGenerator[1106] = 8'hfe;
assign _c_characterGenerator[1107] = 8'h66;
assign _c_characterGenerator[1108] = 8'h62;
assign _c_characterGenerator[1109] = 8'h68;
assign _c_characterGenerator[1110] = 8'h78;
assign _c_characterGenerator[1111] = 8'h68;
assign _c_characterGenerator[1112] = 8'h60;
assign _c_characterGenerator[1113] = 8'h62;
assign _c_characterGenerator[1114] = 8'h66;
assign _c_characterGenerator[1115] = 8'hfe;
assign _c_characterGenerator[1116] = 8'h00;
assign _c_characterGenerator[1117] = 8'h00;
assign _c_characterGenerator[1118] = 8'h00;
assign _c_characterGenerator[1119] = 8'h00;
assign _c_characterGenerator[1120] = 8'h00;
assign _c_characterGenerator[1121] = 8'h00;
assign _c_characterGenerator[1122] = 8'hfe;
assign _c_characterGenerator[1123] = 8'h66;
assign _c_characterGenerator[1124] = 8'h62;
assign _c_characterGenerator[1125] = 8'h68;
assign _c_characterGenerator[1126] = 8'h78;
assign _c_characterGenerator[1127] = 8'h68;
assign _c_characterGenerator[1128] = 8'h60;
assign _c_characterGenerator[1129] = 8'h60;
assign _c_characterGenerator[1130] = 8'h60;
assign _c_characterGenerator[1131] = 8'hf0;
assign _c_characterGenerator[1132] = 8'h00;
assign _c_characterGenerator[1133] = 8'h00;
assign _c_characterGenerator[1134] = 8'h00;
assign _c_characterGenerator[1135] = 8'h00;
assign _c_characterGenerator[1136] = 8'h00;
assign _c_characterGenerator[1137] = 8'h00;
assign _c_characterGenerator[1138] = 8'h3c;
assign _c_characterGenerator[1139] = 8'h66;
assign _c_characterGenerator[1140] = 8'hc2;
assign _c_characterGenerator[1141] = 8'hc0;
assign _c_characterGenerator[1142] = 8'hc0;
assign _c_characterGenerator[1143] = 8'hde;
assign _c_characterGenerator[1144] = 8'hc6;
assign _c_characterGenerator[1145] = 8'hc6;
assign _c_characterGenerator[1146] = 8'h66;
assign _c_characterGenerator[1147] = 8'h3a;
assign _c_characterGenerator[1148] = 8'h00;
assign _c_characterGenerator[1149] = 8'h00;
assign _c_characterGenerator[1150] = 8'h00;
assign _c_characterGenerator[1151] = 8'h00;
assign _c_characterGenerator[1152] = 8'h00;
assign _c_characterGenerator[1153] = 8'h00;
assign _c_characterGenerator[1154] = 8'hc6;
assign _c_characterGenerator[1155] = 8'hc6;
assign _c_characterGenerator[1156] = 8'hc6;
assign _c_characterGenerator[1157] = 8'hc6;
assign _c_characterGenerator[1158] = 8'hfe;
assign _c_characterGenerator[1159] = 8'hc6;
assign _c_characterGenerator[1160] = 8'hc6;
assign _c_characterGenerator[1161] = 8'hc6;
assign _c_characterGenerator[1162] = 8'hc6;
assign _c_characterGenerator[1163] = 8'hc6;
assign _c_characterGenerator[1164] = 8'h00;
assign _c_characterGenerator[1165] = 8'h00;
assign _c_characterGenerator[1166] = 8'h00;
assign _c_characterGenerator[1167] = 8'h00;
assign _c_characterGenerator[1168] = 8'h00;
assign _c_characterGenerator[1169] = 8'h00;
assign _c_characterGenerator[1170] = 8'h3c;
assign _c_characterGenerator[1171] = 8'h18;
assign _c_characterGenerator[1172] = 8'h18;
assign _c_characterGenerator[1173] = 8'h18;
assign _c_characterGenerator[1174] = 8'h18;
assign _c_characterGenerator[1175] = 8'h18;
assign _c_characterGenerator[1176] = 8'h18;
assign _c_characterGenerator[1177] = 8'h18;
assign _c_characterGenerator[1178] = 8'h18;
assign _c_characterGenerator[1179] = 8'h3c;
assign _c_characterGenerator[1180] = 8'h00;
assign _c_characterGenerator[1181] = 8'h00;
assign _c_characterGenerator[1182] = 8'h00;
assign _c_characterGenerator[1183] = 8'h00;
assign _c_characterGenerator[1184] = 8'h00;
assign _c_characterGenerator[1185] = 8'h00;
assign _c_characterGenerator[1186] = 8'h1e;
assign _c_characterGenerator[1187] = 8'h0c;
assign _c_characterGenerator[1188] = 8'h0c;
assign _c_characterGenerator[1189] = 8'h0c;
assign _c_characterGenerator[1190] = 8'h0c;
assign _c_characterGenerator[1191] = 8'h0c;
assign _c_characterGenerator[1192] = 8'hcc;
assign _c_characterGenerator[1193] = 8'hcc;
assign _c_characterGenerator[1194] = 8'hcc;
assign _c_characterGenerator[1195] = 8'h78;
assign _c_characterGenerator[1196] = 8'h00;
assign _c_characterGenerator[1197] = 8'h00;
assign _c_characterGenerator[1198] = 8'h00;
assign _c_characterGenerator[1199] = 8'h00;
assign _c_characterGenerator[1200] = 8'h00;
assign _c_characterGenerator[1201] = 8'h00;
assign _c_characterGenerator[1202] = 8'he6;
assign _c_characterGenerator[1203] = 8'h66;
assign _c_characterGenerator[1204] = 8'h66;
assign _c_characterGenerator[1205] = 8'h6c;
assign _c_characterGenerator[1206] = 8'h78;
assign _c_characterGenerator[1207] = 8'h78;
assign _c_characterGenerator[1208] = 8'h6c;
assign _c_characterGenerator[1209] = 8'h66;
assign _c_characterGenerator[1210] = 8'h66;
assign _c_characterGenerator[1211] = 8'he6;
assign _c_characterGenerator[1212] = 8'h00;
assign _c_characterGenerator[1213] = 8'h00;
assign _c_characterGenerator[1214] = 8'h00;
assign _c_characterGenerator[1215] = 8'h00;
assign _c_characterGenerator[1216] = 8'h00;
assign _c_characterGenerator[1217] = 8'h00;
assign _c_characterGenerator[1218] = 8'hf0;
assign _c_characterGenerator[1219] = 8'h60;
assign _c_characterGenerator[1220] = 8'h60;
assign _c_characterGenerator[1221] = 8'h60;
assign _c_characterGenerator[1222] = 8'h60;
assign _c_characterGenerator[1223] = 8'h60;
assign _c_characterGenerator[1224] = 8'h60;
assign _c_characterGenerator[1225] = 8'h62;
assign _c_characterGenerator[1226] = 8'h66;
assign _c_characterGenerator[1227] = 8'hfe;
assign _c_characterGenerator[1228] = 8'h00;
assign _c_characterGenerator[1229] = 8'h00;
assign _c_characterGenerator[1230] = 8'h00;
assign _c_characterGenerator[1231] = 8'h00;
assign _c_characterGenerator[1232] = 8'h00;
assign _c_characterGenerator[1233] = 8'h00;
assign _c_characterGenerator[1234] = 8'hc6;
assign _c_characterGenerator[1235] = 8'hee;
assign _c_characterGenerator[1236] = 8'hfe;
assign _c_characterGenerator[1237] = 8'hfe;
assign _c_characterGenerator[1238] = 8'hd6;
assign _c_characterGenerator[1239] = 8'hc6;
assign _c_characterGenerator[1240] = 8'hc6;
assign _c_characterGenerator[1241] = 8'hc6;
assign _c_characterGenerator[1242] = 8'hc6;
assign _c_characterGenerator[1243] = 8'hc6;
assign _c_characterGenerator[1244] = 8'h00;
assign _c_characterGenerator[1245] = 8'h00;
assign _c_characterGenerator[1246] = 8'h00;
assign _c_characterGenerator[1247] = 8'h00;
assign _c_characterGenerator[1248] = 8'h00;
assign _c_characterGenerator[1249] = 8'h00;
assign _c_characterGenerator[1250] = 8'hc6;
assign _c_characterGenerator[1251] = 8'he6;
assign _c_characterGenerator[1252] = 8'hf6;
assign _c_characterGenerator[1253] = 8'hfe;
assign _c_characterGenerator[1254] = 8'hde;
assign _c_characterGenerator[1255] = 8'hce;
assign _c_characterGenerator[1256] = 8'hc6;
assign _c_characterGenerator[1257] = 8'hc6;
assign _c_characterGenerator[1258] = 8'hc6;
assign _c_characterGenerator[1259] = 8'hc6;
assign _c_characterGenerator[1260] = 8'h00;
assign _c_characterGenerator[1261] = 8'h00;
assign _c_characterGenerator[1262] = 8'h00;
assign _c_characterGenerator[1263] = 8'h00;
assign _c_characterGenerator[1264] = 8'h00;
assign _c_characterGenerator[1265] = 8'h00;
assign _c_characterGenerator[1266] = 8'h7c;
assign _c_characterGenerator[1267] = 8'hc6;
assign _c_characterGenerator[1268] = 8'hc6;
assign _c_characterGenerator[1269] = 8'hc6;
assign _c_characterGenerator[1270] = 8'hc6;
assign _c_characterGenerator[1271] = 8'hc6;
assign _c_characterGenerator[1272] = 8'hc6;
assign _c_characterGenerator[1273] = 8'hc6;
assign _c_characterGenerator[1274] = 8'hc6;
assign _c_characterGenerator[1275] = 8'h7c;
assign _c_characterGenerator[1276] = 8'h00;
assign _c_characterGenerator[1277] = 8'h00;
assign _c_characterGenerator[1278] = 8'h00;
assign _c_characterGenerator[1279] = 8'h00;
assign _c_characterGenerator[1280] = 8'h00;
assign _c_characterGenerator[1281] = 8'h00;
assign _c_characterGenerator[1282] = 8'hfc;
assign _c_characterGenerator[1283] = 8'h66;
assign _c_characterGenerator[1284] = 8'h66;
assign _c_characterGenerator[1285] = 8'h66;
assign _c_characterGenerator[1286] = 8'h7c;
assign _c_characterGenerator[1287] = 8'h60;
assign _c_characterGenerator[1288] = 8'h60;
assign _c_characterGenerator[1289] = 8'h60;
assign _c_characterGenerator[1290] = 8'h60;
assign _c_characterGenerator[1291] = 8'hf0;
assign _c_characterGenerator[1292] = 8'h00;
assign _c_characterGenerator[1293] = 8'h00;
assign _c_characterGenerator[1294] = 8'h00;
assign _c_characterGenerator[1295] = 8'h00;
assign _c_characterGenerator[1296] = 8'h00;
assign _c_characterGenerator[1297] = 8'h00;
assign _c_characterGenerator[1298] = 8'h7c;
assign _c_characterGenerator[1299] = 8'hc6;
assign _c_characterGenerator[1300] = 8'hc6;
assign _c_characterGenerator[1301] = 8'hc6;
assign _c_characterGenerator[1302] = 8'hc6;
assign _c_characterGenerator[1303] = 8'hc6;
assign _c_characterGenerator[1304] = 8'hc6;
assign _c_characterGenerator[1305] = 8'hd6;
assign _c_characterGenerator[1306] = 8'hde;
assign _c_characterGenerator[1307] = 8'h7c;
assign _c_characterGenerator[1308] = 8'h0c;
assign _c_characterGenerator[1309] = 8'h0e;
assign _c_characterGenerator[1310] = 8'h00;
assign _c_characterGenerator[1311] = 8'h00;
assign _c_characterGenerator[1312] = 8'h00;
assign _c_characterGenerator[1313] = 8'h00;
assign _c_characterGenerator[1314] = 8'hfc;
assign _c_characterGenerator[1315] = 8'h66;
assign _c_characterGenerator[1316] = 8'h66;
assign _c_characterGenerator[1317] = 8'h66;
assign _c_characterGenerator[1318] = 8'h7c;
assign _c_characterGenerator[1319] = 8'h6c;
assign _c_characterGenerator[1320] = 8'h66;
assign _c_characterGenerator[1321] = 8'h66;
assign _c_characterGenerator[1322] = 8'h66;
assign _c_characterGenerator[1323] = 8'he6;
assign _c_characterGenerator[1324] = 8'h00;
assign _c_characterGenerator[1325] = 8'h00;
assign _c_characterGenerator[1326] = 8'h00;
assign _c_characterGenerator[1327] = 8'h00;
assign _c_characterGenerator[1328] = 8'h00;
assign _c_characterGenerator[1329] = 8'h00;
assign _c_characterGenerator[1330] = 8'h7c;
assign _c_characterGenerator[1331] = 8'hc6;
assign _c_characterGenerator[1332] = 8'hc6;
assign _c_characterGenerator[1333] = 8'h60;
assign _c_characterGenerator[1334] = 8'h38;
assign _c_characterGenerator[1335] = 8'h0c;
assign _c_characterGenerator[1336] = 8'h06;
assign _c_characterGenerator[1337] = 8'hc6;
assign _c_characterGenerator[1338] = 8'hc6;
assign _c_characterGenerator[1339] = 8'h7c;
assign _c_characterGenerator[1340] = 8'h00;
assign _c_characterGenerator[1341] = 8'h00;
assign _c_characterGenerator[1342] = 8'h00;
assign _c_characterGenerator[1343] = 8'h00;
assign _c_characterGenerator[1344] = 8'h00;
assign _c_characterGenerator[1345] = 8'h00;
assign _c_characterGenerator[1346] = 8'h7e;
assign _c_characterGenerator[1347] = 8'h7e;
assign _c_characterGenerator[1348] = 8'h5a;
assign _c_characterGenerator[1349] = 8'h18;
assign _c_characterGenerator[1350] = 8'h18;
assign _c_characterGenerator[1351] = 8'h18;
assign _c_characterGenerator[1352] = 8'h18;
assign _c_characterGenerator[1353] = 8'h18;
assign _c_characterGenerator[1354] = 8'h18;
assign _c_characterGenerator[1355] = 8'h3c;
assign _c_characterGenerator[1356] = 8'h00;
assign _c_characterGenerator[1357] = 8'h00;
assign _c_characterGenerator[1358] = 8'h00;
assign _c_characterGenerator[1359] = 8'h00;
assign _c_characterGenerator[1360] = 8'h00;
assign _c_characterGenerator[1361] = 8'h00;
assign _c_characterGenerator[1362] = 8'hc6;
assign _c_characterGenerator[1363] = 8'hc6;
assign _c_characterGenerator[1364] = 8'hc6;
assign _c_characterGenerator[1365] = 8'hc6;
assign _c_characterGenerator[1366] = 8'hc6;
assign _c_characterGenerator[1367] = 8'hc6;
assign _c_characterGenerator[1368] = 8'hc6;
assign _c_characterGenerator[1369] = 8'hc6;
assign _c_characterGenerator[1370] = 8'hc6;
assign _c_characterGenerator[1371] = 8'h7c;
assign _c_characterGenerator[1372] = 8'h00;
assign _c_characterGenerator[1373] = 8'h00;
assign _c_characterGenerator[1374] = 8'h00;
assign _c_characterGenerator[1375] = 8'h00;
assign _c_characterGenerator[1376] = 8'h00;
assign _c_characterGenerator[1377] = 8'h00;
assign _c_characterGenerator[1378] = 8'hc6;
assign _c_characterGenerator[1379] = 8'hc6;
assign _c_characterGenerator[1380] = 8'hc6;
assign _c_characterGenerator[1381] = 8'hc6;
assign _c_characterGenerator[1382] = 8'hc6;
assign _c_characterGenerator[1383] = 8'hc6;
assign _c_characterGenerator[1384] = 8'hc6;
assign _c_characterGenerator[1385] = 8'h6c;
assign _c_characterGenerator[1386] = 8'h38;
assign _c_characterGenerator[1387] = 8'h10;
assign _c_characterGenerator[1388] = 8'h00;
assign _c_characterGenerator[1389] = 8'h00;
assign _c_characterGenerator[1390] = 8'h00;
assign _c_characterGenerator[1391] = 8'h00;
assign _c_characterGenerator[1392] = 8'h00;
assign _c_characterGenerator[1393] = 8'h00;
assign _c_characterGenerator[1394] = 8'hc6;
assign _c_characterGenerator[1395] = 8'hc6;
assign _c_characterGenerator[1396] = 8'hc6;
assign _c_characterGenerator[1397] = 8'hc6;
assign _c_characterGenerator[1398] = 8'hd6;
assign _c_characterGenerator[1399] = 8'hd6;
assign _c_characterGenerator[1400] = 8'hd6;
assign _c_characterGenerator[1401] = 8'hfe;
assign _c_characterGenerator[1402] = 8'hee;
assign _c_characterGenerator[1403] = 8'h6c;
assign _c_characterGenerator[1404] = 8'h00;
assign _c_characterGenerator[1405] = 8'h00;
assign _c_characterGenerator[1406] = 8'h00;
assign _c_characterGenerator[1407] = 8'h00;
assign _c_characterGenerator[1408] = 8'h00;
assign _c_characterGenerator[1409] = 8'h00;
assign _c_characterGenerator[1410] = 8'hc6;
assign _c_characterGenerator[1411] = 8'hc6;
assign _c_characterGenerator[1412] = 8'h6c;
assign _c_characterGenerator[1413] = 8'h7c;
assign _c_characterGenerator[1414] = 8'h38;
assign _c_characterGenerator[1415] = 8'h38;
assign _c_characterGenerator[1416] = 8'h7c;
assign _c_characterGenerator[1417] = 8'h6c;
assign _c_characterGenerator[1418] = 8'hc6;
assign _c_characterGenerator[1419] = 8'hc6;
assign _c_characterGenerator[1420] = 8'h00;
assign _c_characterGenerator[1421] = 8'h00;
assign _c_characterGenerator[1422] = 8'h00;
assign _c_characterGenerator[1423] = 8'h00;
assign _c_characterGenerator[1424] = 8'h00;
assign _c_characterGenerator[1425] = 8'h00;
assign _c_characterGenerator[1426] = 8'h66;
assign _c_characterGenerator[1427] = 8'h66;
assign _c_characterGenerator[1428] = 8'h66;
assign _c_characterGenerator[1429] = 8'h66;
assign _c_characterGenerator[1430] = 8'h3c;
assign _c_characterGenerator[1431] = 8'h18;
assign _c_characterGenerator[1432] = 8'h18;
assign _c_characterGenerator[1433] = 8'h18;
assign _c_characterGenerator[1434] = 8'h18;
assign _c_characterGenerator[1435] = 8'h3c;
assign _c_characterGenerator[1436] = 8'h00;
assign _c_characterGenerator[1437] = 8'h00;
assign _c_characterGenerator[1438] = 8'h00;
assign _c_characterGenerator[1439] = 8'h00;
assign _c_characterGenerator[1440] = 8'h00;
assign _c_characterGenerator[1441] = 8'h00;
assign _c_characterGenerator[1442] = 8'hfe;
assign _c_characterGenerator[1443] = 8'hc6;
assign _c_characterGenerator[1444] = 8'h86;
assign _c_characterGenerator[1445] = 8'h0c;
assign _c_characterGenerator[1446] = 8'h18;
assign _c_characterGenerator[1447] = 8'h30;
assign _c_characterGenerator[1448] = 8'h60;
assign _c_characterGenerator[1449] = 8'hc2;
assign _c_characterGenerator[1450] = 8'hc6;
assign _c_characterGenerator[1451] = 8'hfe;
assign _c_characterGenerator[1452] = 8'h00;
assign _c_characterGenerator[1453] = 8'h00;
assign _c_characterGenerator[1454] = 8'h00;
assign _c_characterGenerator[1455] = 8'h00;
assign _c_characterGenerator[1456] = 8'h00;
assign _c_characterGenerator[1457] = 8'h00;
assign _c_characterGenerator[1458] = 8'h3c;
assign _c_characterGenerator[1459] = 8'h30;
assign _c_characterGenerator[1460] = 8'h30;
assign _c_characterGenerator[1461] = 8'h30;
assign _c_characterGenerator[1462] = 8'h30;
assign _c_characterGenerator[1463] = 8'h30;
assign _c_characterGenerator[1464] = 8'h30;
assign _c_characterGenerator[1465] = 8'h30;
assign _c_characterGenerator[1466] = 8'h30;
assign _c_characterGenerator[1467] = 8'h3c;
assign _c_characterGenerator[1468] = 8'h00;
assign _c_characterGenerator[1469] = 8'h00;
assign _c_characterGenerator[1470] = 8'h00;
assign _c_characterGenerator[1471] = 8'h00;
assign _c_characterGenerator[1472] = 8'h00;
assign _c_characterGenerator[1473] = 8'h00;
assign _c_characterGenerator[1474] = 8'h00;
assign _c_characterGenerator[1475] = 8'h80;
assign _c_characterGenerator[1476] = 8'hc0;
assign _c_characterGenerator[1477] = 8'he0;
assign _c_characterGenerator[1478] = 8'h70;
assign _c_characterGenerator[1479] = 8'h38;
assign _c_characterGenerator[1480] = 8'h1c;
assign _c_characterGenerator[1481] = 8'h0e;
assign _c_characterGenerator[1482] = 8'h06;
assign _c_characterGenerator[1483] = 8'h02;
assign _c_characterGenerator[1484] = 8'h00;
assign _c_characterGenerator[1485] = 8'h00;
assign _c_characterGenerator[1486] = 8'h00;
assign _c_characterGenerator[1487] = 8'h00;
assign _c_characterGenerator[1488] = 8'h00;
assign _c_characterGenerator[1489] = 8'h00;
assign _c_characterGenerator[1490] = 8'h3c;
assign _c_characterGenerator[1491] = 8'h0c;
assign _c_characterGenerator[1492] = 8'h0c;
assign _c_characterGenerator[1493] = 8'h0c;
assign _c_characterGenerator[1494] = 8'h0c;
assign _c_characterGenerator[1495] = 8'h0c;
assign _c_characterGenerator[1496] = 8'h0c;
assign _c_characterGenerator[1497] = 8'h0c;
assign _c_characterGenerator[1498] = 8'h0c;
assign _c_characterGenerator[1499] = 8'h3c;
assign _c_characterGenerator[1500] = 8'h00;
assign _c_characterGenerator[1501] = 8'h00;
assign _c_characterGenerator[1502] = 8'h00;
assign _c_characterGenerator[1503] = 8'h00;
assign _c_characterGenerator[1504] = 8'h10;
assign _c_characterGenerator[1505] = 8'h38;
assign _c_characterGenerator[1506] = 8'h6c;
assign _c_characterGenerator[1507] = 8'hc6;
assign _c_characterGenerator[1508] = 8'h00;
assign _c_characterGenerator[1509] = 8'h00;
assign _c_characterGenerator[1510] = 8'h00;
assign _c_characterGenerator[1511] = 8'h00;
assign _c_characterGenerator[1512] = 8'h00;
assign _c_characterGenerator[1513] = 8'h00;
assign _c_characterGenerator[1514] = 8'h00;
assign _c_characterGenerator[1515] = 8'h00;
assign _c_characterGenerator[1516] = 8'h00;
assign _c_characterGenerator[1517] = 8'h00;
assign _c_characterGenerator[1518] = 8'h00;
assign _c_characterGenerator[1519] = 8'h00;
assign _c_characterGenerator[1520] = 8'h00;
assign _c_characterGenerator[1521] = 8'h00;
assign _c_characterGenerator[1522] = 8'h00;
assign _c_characterGenerator[1523] = 8'h00;
assign _c_characterGenerator[1524] = 8'h00;
assign _c_characterGenerator[1525] = 8'h00;
assign _c_characterGenerator[1526] = 8'h00;
assign _c_characterGenerator[1527] = 8'h00;
assign _c_characterGenerator[1528] = 8'h00;
assign _c_characterGenerator[1529] = 8'h00;
assign _c_characterGenerator[1530] = 8'h00;
assign _c_characterGenerator[1531] = 8'h00;
assign _c_characterGenerator[1532] = 8'h00;
assign _c_characterGenerator[1533] = 8'hff;
assign _c_characterGenerator[1534] = 8'h00;
assign _c_characterGenerator[1535] = 8'h00;
assign _c_characterGenerator[1536] = 8'h30;
assign _c_characterGenerator[1537] = 8'h30;
assign _c_characterGenerator[1538] = 8'h18;
assign _c_characterGenerator[1539] = 8'h00;
assign _c_characterGenerator[1540] = 8'h00;
assign _c_characterGenerator[1541] = 8'h00;
assign _c_characterGenerator[1542] = 8'h00;
assign _c_characterGenerator[1543] = 8'h00;
assign _c_characterGenerator[1544] = 8'h00;
assign _c_characterGenerator[1545] = 8'h00;
assign _c_characterGenerator[1546] = 8'h00;
assign _c_characterGenerator[1547] = 8'h00;
assign _c_characterGenerator[1548] = 8'h00;
assign _c_characterGenerator[1549] = 8'h00;
assign _c_characterGenerator[1550] = 8'h00;
assign _c_characterGenerator[1551] = 8'h00;
assign _c_characterGenerator[1552] = 8'h00;
assign _c_characterGenerator[1553] = 8'h00;
assign _c_characterGenerator[1554] = 8'h00;
assign _c_characterGenerator[1555] = 8'h00;
assign _c_characterGenerator[1556] = 8'h00;
assign _c_characterGenerator[1557] = 8'h78;
assign _c_characterGenerator[1558] = 8'h0c;
assign _c_characterGenerator[1559] = 8'h7c;
assign _c_characterGenerator[1560] = 8'hcc;
assign _c_characterGenerator[1561] = 8'hcc;
assign _c_characterGenerator[1562] = 8'hcc;
assign _c_characterGenerator[1563] = 8'h76;
assign _c_characterGenerator[1564] = 8'h00;
assign _c_characterGenerator[1565] = 8'h00;
assign _c_characterGenerator[1566] = 8'h00;
assign _c_characterGenerator[1567] = 8'h00;
assign _c_characterGenerator[1568] = 8'h00;
assign _c_characterGenerator[1569] = 8'h00;
assign _c_characterGenerator[1570] = 8'he0;
assign _c_characterGenerator[1571] = 8'h60;
assign _c_characterGenerator[1572] = 8'h60;
assign _c_characterGenerator[1573] = 8'h78;
assign _c_characterGenerator[1574] = 8'h6c;
assign _c_characterGenerator[1575] = 8'h66;
assign _c_characterGenerator[1576] = 8'h66;
assign _c_characterGenerator[1577] = 8'h66;
assign _c_characterGenerator[1578] = 8'h66;
assign _c_characterGenerator[1579] = 8'h7c;
assign _c_characterGenerator[1580] = 8'h00;
assign _c_characterGenerator[1581] = 8'h00;
assign _c_characterGenerator[1582] = 8'h00;
assign _c_characterGenerator[1583] = 8'h00;
assign _c_characterGenerator[1584] = 8'h00;
assign _c_characterGenerator[1585] = 8'h00;
assign _c_characterGenerator[1586] = 8'h00;
assign _c_characterGenerator[1587] = 8'h00;
assign _c_characterGenerator[1588] = 8'h00;
assign _c_characterGenerator[1589] = 8'h7c;
assign _c_characterGenerator[1590] = 8'hc6;
assign _c_characterGenerator[1591] = 8'hc0;
assign _c_characterGenerator[1592] = 8'hc0;
assign _c_characterGenerator[1593] = 8'hc0;
assign _c_characterGenerator[1594] = 8'hc6;
assign _c_characterGenerator[1595] = 8'h7c;
assign _c_characterGenerator[1596] = 8'h00;
assign _c_characterGenerator[1597] = 8'h00;
assign _c_characterGenerator[1598] = 8'h00;
assign _c_characterGenerator[1599] = 8'h00;
assign _c_characterGenerator[1600] = 8'h00;
assign _c_characterGenerator[1601] = 8'h00;
assign _c_characterGenerator[1602] = 8'h1c;
assign _c_characterGenerator[1603] = 8'h0c;
assign _c_characterGenerator[1604] = 8'h0c;
assign _c_characterGenerator[1605] = 8'h3c;
assign _c_characterGenerator[1606] = 8'h6c;
assign _c_characterGenerator[1607] = 8'hcc;
assign _c_characterGenerator[1608] = 8'hcc;
assign _c_characterGenerator[1609] = 8'hcc;
assign _c_characterGenerator[1610] = 8'hcc;
assign _c_characterGenerator[1611] = 8'h76;
assign _c_characterGenerator[1612] = 8'h00;
assign _c_characterGenerator[1613] = 8'h00;
assign _c_characterGenerator[1614] = 8'h00;
assign _c_characterGenerator[1615] = 8'h00;
assign _c_characterGenerator[1616] = 8'h00;
assign _c_characterGenerator[1617] = 8'h00;
assign _c_characterGenerator[1618] = 8'h00;
assign _c_characterGenerator[1619] = 8'h00;
assign _c_characterGenerator[1620] = 8'h00;
assign _c_characterGenerator[1621] = 8'h7c;
assign _c_characterGenerator[1622] = 8'hc6;
assign _c_characterGenerator[1623] = 8'hfe;
assign _c_characterGenerator[1624] = 8'hc0;
assign _c_characterGenerator[1625] = 8'hc0;
assign _c_characterGenerator[1626] = 8'hc6;
assign _c_characterGenerator[1627] = 8'h7c;
assign _c_characterGenerator[1628] = 8'h00;
assign _c_characterGenerator[1629] = 8'h00;
assign _c_characterGenerator[1630] = 8'h00;
assign _c_characterGenerator[1631] = 8'h00;
assign _c_characterGenerator[1632] = 8'h00;
assign _c_characterGenerator[1633] = 8'h00;
assign _c_characterGenerator[1634] = 8'h38;
assign _c_characterGenerator[1635] = 8'h6c;
assign _c_characterGenerator[1636] = 8'h64;
assign _c_characterGenerator[1637] = 8'h60;
assign _c_characterGenerator[1638] = 8'hf0;
assign _c_characterGenerator[1639] = 8'h60;
assign _c_characterGenerator[1640] = 8'h60;
assign _c_characterGenerator[1641] = 8'h60;
assign _c_characterGenerator[1642] = 8'h60;
assign _c_characterGenerator[1643] = 8'hf0;
assign _c_characterGenerator[1644] = 8'h00;
assign _c_characterGenerator[1645] = 8'h00;
assign _c_characterGenerator[1646] = 8'h00;
assign _c_characterGenerator[1647] = 8'h00;
assign _c_characterGenerator[1648] = 8'h00;
assign _c_characterGenerator[1649] = 8'h00;
assign _c_characterGenerator[1650] = 8'h00;
assign _c_characterGenerator[1651] = 8'h00;
assign _c_characterGenerator[1652] = 8'h00;
assign _c_characterGenerator[1653] = 8'h76;
assign _c_characterGenerator[1654] = 8'hcc;
assign _c_characterGenerator[1655] = 8'hcc;
assign _c_characterGenerator[1656] = 8'hcc;
assign _c_characterGenerator[1657] = 8'hcc;
assign _c_characterGenerator[1658] = 8'hcc;
assign _c_characterGenerator[1659] = 8'h7c;
assign _c_characterGenerator[1660] = 8'h0c;
assign _c_characterGenerator[1661] = 8'hcc;
assign _c_characterGenerator[1662] = 8'h78;
assign _c_characterGenerator[1663] = 8'h00;
assign _c_characterGenerator[1664] = 8'h00;
assign _c_characterGenerator[1665] = 8'h00;
assign _c_characterGenerator[1666] = 8'he0;
assign _c_characterGenerator[1667] = 8'h60;
assign _c_characterGenerator[1668] = 8'h60;
assign _c_characterGenerator[1669] = 8'h6c;
assign _c_characterGenerator[1670] = 8'h76;
assign _c_characterGenerator[1671] = 8'h66;
assign _c_characterGenerator[1672] = 8'h66;
assign _c_characterGenerator[1673] = 8'h66;
assign _c_characterGenerator[1674] = 8'h66;
assign _c_characterGenerator[1675] = 8'he6;
assign _c_characterGenerator[1676] = 8'h00;
assign _c_characterGenerator[1677] = 8'h00;
assign _c_characterGenerator[1678] = 8'h00;
assign _c_characterGenerator[1679] = 8'h00;
assign _c_characterGenerator[1680] = 8'h00;
assign _c_characterGenerator[1681] = 8'h00;
assign _c_characterGenerator[1682] = 8'h18;
assign _c_characterGenerator[1683] = 8'h18;
assign _c_characterGenerator[1684] = 8'h00;
assign _c_characterGenerator[1685] = 8'h38;
assign _c_characterGenerator[1686] = 8'h18;
assign _c_characterGenerator[1687] = 8'h18;
assign _c_characterGenerator[1688] = 8'h18;
assign _c_characterGenerator[1689] = 8'h18;
assign _c_characterGenerator[1690] = 8'h18;
assign _c_characterGenerator[1691] = 8'h3c;
assign _c_characterGenerator[1692] = 8'h00;
assign _c_characterGenerator[1693] = 8'h00;
assign _c_characterGenerator[1694] = 8'h00;
assign _c_characterGenerator[1695] = 8'h00;
assign _c_characterGenerator[1696] = 8'h00;
assign _c_characterGenerator[1697] = 8'h00;
assign _c_characterGenerator[1698] = 8'h06;
assign _c_characterGenerator[1699] = 8'h06;
assign _c_characterGenerator[1700] = 8'h00;
assign _c_characterGenerator[1701] = 8'h0e;
assign _c_characterGenerator[1702] = 8'h06;
assign _c_characterGenerator[1703] = 8'h06;
assign _c_characterGenerator[1704] = 8'h06;
assign _c_characterGenerator[1705] = 8'h06;
assign _c_characterGenerator[1706] = 8'h06;
assign _c_characterGenerator[1707] = 8'h06;
assign _c_characterGenerator[1708] = 8'h66;
assign _c_characterGenerator[1709] = 8'h66;
assign _c_characterGenerator[1710] = 8'h3c;
assign _c_characterGenerator[1711] = 8'h00;
assign _c_characterGenerator[1712] = 8'h00;
assign _c_characterGenerator[1713] = 8'h00;
assign _c_characterGenerator[1714] = 8'he0;
assign _c_characterGenerator[1715] = 8'h60;
assign _c_characterGenerator[1716] = 8'h60;
assign _c_characterGenerator[1717] = 8'h66;
assign _c_characterGenerator[1718] = 8'h6c;
assign _c_characterGenerator[1719] = 8'h78;
assign _c_characterGenerator[1720] = 8'h78;
assign _c_characterGenerator[1721] = 8'h6c;
assign _c_characterGenerator[1722] = 8'h66;
assign _c_characterGenerator[1723] = 8'he6;
assign _c_characterGenerator[1724] = 8'h00;
assign _c_characterGenerator[1725] = 8'h00;
assign _c_characterGenerator[1726] = 8'h00;
assign _c_characterGenerator[1727] = 8'h00;
assign _c_characterGenerator[1728] = 8'h00;
assign _c_characterGenerator[1729] = 8'h00;
assign _c_characterGenerator[1730] = 8'h38;
assign _c_characterGenerator[1731] = 8'h18;
assign _c_characterGenerator[1732] = 8'h18;
assign _c_characterGenerator[1733] = 8'h18;
assign _c_characterGenerator[1734] = 8'h18;
assign _c_characterGenerator[1735] = 8'h18;
assign _c_characterGenerator[1736] = 8'h18;
assign _c_characterGenerator[1737] = 8'h18;
assign _c_characterGenerator[1738] = 8'h18;
assign _c_characterGenerator[1739] = 8'h3c;
assign _c_characterGenerator[1740] = 8'h00;
assign _c_characterGenerator[1741] = 8'h00;
assign _c_characterGenerator[1742] = 8'h00;
assign _c_characterGenerator[1743] = 8'h00;
assign _c_characterGenerator[1744] = 8'h00;
assign _c_characterGenerator[1745] = 8'h00;
assign _c_characterGenerator[1746] = 8'h00;
assign _c_characterGenerator[1747] = 8'h00;
assign _c_characterGenerator[1748] = 8'h00;
assign _c_characterGenerator[1749] = 8'hec;
assign _c_characterGenerator[1750] = 8'hfe;
assign _c_characterGenerator[1751] = 8'hd6;
assign _c_characterGenerator[1752] = 8'hd6;
assign _c_characterGenerator[1753] = 8'hd6;
assign _c_characterGenerator[1754] = 8'hd6;
assign _c_characterGenerator[1755] = 8'hc6;
assign _c_characterGenerator[1756] = 8'h00;
assign _c_characterGenerator[1757] = 8'h00;
assign _c_characterGenerator[1758] = 8'h00;
assign _c_characterGenerator[1759] = 8'h00;
assign _c_characterGenerator[1760] = 8'h00;
assign _c_characterGenerator[1761] = 8'h00;
assign _c_characterGenerator[1762] = 8'h00;
assign _c_characterGenerator[1763] = 8'h00;
assign _c_characterGenerator[1764] = 8'h00;
assign _c_characterGenerator[1765] = 8'hdc;
assign _c_characterGenerator[1766] = 8'h66;
assign _c_characterGenerator[1767] = 8'h66;
assign _c_characterGenerator[1768] = 8'h66;
assign _c_characterGenerator[1769] = 8'h66;
assign _c_characterGenerator[1770] = 8'h66;
assign _c_characterGenerator[1771] = 8'h66;
assign _c_characterGenerator[1772] = 8'h00;
assign _c_characterGenerator[1773] = 8'h00;
assign _c_characterGenerator[1774] = 8'h00;
assign _c_characterGenerator[1775] = 8'h00;
assign _c_characterGenerator[1776] = 8'h00;
assign _c_characterGenerator[1777] = 8'h00;
assign _c_characterGenerator[1778] = 8'h00;
assign _c_characterGenerator[1779] = 8'h00;
assign _c_characterGenerator[1780] = 8'h00;
assign _c_characterGenerator[1781] = 8'h7c;
assign _c_characterGenerator[1782] = 8'hc6;
assign _c_characterGenerator[1783] = 8'hc6;
assign _c_characterGenerator[1784] = 8'hc6;
assign _c_characterGenerator[1785] = 8'hc6;
assign _c_characterGenerator[1786] = 8'hc6;
assign _c_characterGenerator[1787] = 8'h7c;
assign _c_characterGenerator[1788] = 8'h00;
assign _c_characterGenerator[1789] = 8'h00;
assign _c_characterGenerator[1790] = 8'h00;
assign _c_characterGenerator[1791] = 8'h00;
assign _c_characterGenerator[1792] = 8'h00;
assign _c_characterGenerator[1793] = 8'h00;
assign _c_characterGenerator[1794] = 8'h00;
assign _c_characterGenerator[1795] = 8'h00;
assign _c_characterGenerator[1796] = 8'h00;
assign _c_characterGenerator[1797] = 8'hdc;
assign _c_characterGenerator[1798] = 8'h66;
assign _c_characterGenerator[1799] = 8'h66;
assign _c_characterGenerator[1800] = 8'h66;
assign _c_characterGenerator[1801] = 8'h66;
assign _c_characterGenerator[1802] = 8'h66;
assign _c_characterGenerator[1803] = 8'h7c;
assign _c_characterGenerator[1804] = 8'h60;
assign _c_characterGenerator[1805] = 8'h60;
assign _c_characterGenerator[1806] = 8'hf0;
assign _c_characterGenerator[1807] = 8'h00;
assign _c_characterGenerator[1808] = 8'h00;
assign _c_characterGenerator[1809] = 8'h00;
assign _c_characterGenerator[1810] = 8'h00;
assign _c_characterGenerator[1811] = 8'h00;
assign _c_characterGenerator[1812] = 8'h00;
assign _c_characterGenerator[1813] = 8'h76;
assign _c_characterGenerator[1814] = 8'hcc;
assign _c_characterGenerator[1815] = 8'hcc;
assign _c_characterGenerator[1816] = 8'hcc;
assign _c_characterGenerator[1817] = 8'hcc;
assign _c_characterGenerator[1818] = 8'hcc;
assign _c_characterGenerator[1819] = 8'h7c;
assign _c_characterGenerator[1820] = 8'h0c;
assign _c_characterGenerator[1821] = 8'h0c;
assign _c_characterGenerator[1822] = 8'h1e;
assign _c_characterGenerator[1823] = 8'h00;
assign _c_characterGenerator[1824] = 8'h00;
assign _c_characterGenerator[1825] = 8'h00;
assign _c_characterGenerator[1826] = 8'h00;
assign _c_characterGenerator[1827] = 8'h00;
assign _c_characterGenerator[1828] = 8'h00;
assign _c_characterGenerator[1829] = 8'hdc;
assign _c_characterGenerator[1830] = 8'h76;
assign _c_characterGenerator[1831] = 8'h66;
assign _c_characterGenerator[1832] = 8'h60;
assign _c_characterGenerator[1833] = 8'h60;
assign _c_characterGenerator[1834] = 8'h60;
assign _c_characterGenerator[1835] = 8'hf0;
assign _c_characterGenerator[1836] = 8'h00;
assign _c_characterGenerator[1837] = 8'h00;
assign _c_characterGenerator[1838] = 8'h00;
assign _c_characterGenerator[1839] = 8'h00;
assign _c_characterGenerator[1840] = 8'h00;
assign _c_characterGenerator[1841] = 8'h00;
assign _c_characterGenerator[1842] = 8'h00;
assign _c_characterGenerator[1843] = 8'h00;
assign _c_characterGenerator[1844] = 8'h00;
assign _c_characterGenerator[1845] = 8'h7c;
assign _c_characterGenerator[1846] = 8'hc6;
assign _c_characterGenerator[1847] = 8'h60;
assign _c_characterGenerator[1848] = 8'h38;
assign _c_characterGenerator[1849] = 8'h0c;
assign _c_characterGenerator[1850] = 8'hc6;
assign _c_characterGenerator[1851] = 8'h7c;
assign _c_characterGenerator[1852] = 8'h00;
assign _c_characterGenerator[1853] = 8'h00;
assign _c_characterGenerator[1854] = 8'h00;
assign _c_characterGenerator[1855] = 8'h00;
assign _c_characterGenerator[1856] = 8'h00;
assign _c_characterGenerator[1857] = 8'h00;
assign _c_characterGenerator[1858] = 8'h10;
assign _c_characterGenerator[1859] = 8'h30;
assign _c_characterGenerator[1860] = 8'h30;
assign _c_characterGenerator[1861] = 8'hfc;
assign _c_characterGenerator[1862] = 8'h30;
assign _c_characterGenerator[1863] = 8'h30;
assign _c_characterGenerator[1864] = 8'h30;
assign _c_characterGenerator[1865] = 8'h30;
assign _c_characterGenerator[1866] = 8'h36;
assign _c_characterGenerator[1867] = 8'h1c;
assign _c_characterGenerator[1868] = 8'h00;
assign _c_characterGenerator[1869] = 8'h00;
assign _c_characterGenerator[1870] = 8'h00;
assign _c_characterGenerator[1871] = 8'h00;
assign _c_characterGenerator[1872] = 8'h00;
assign _c_characterGenerator[1873] = 8'h00;
assign _c_characterGenerator[1874] = 8'h00;
assign _c_characterGenerator[1875] = 8'h00;
assign _c_characterGenerator[1876] = 8'h00;
assign _c_characterGenerator[1877] = 8'hcc;
assign _c_characterGenerator[1878] = 8'hcc;
assign _c_characterGenerator[1879] = 8'hcc;
assign _c_characterGenerator[1880] = 8'hcc;
assign _c_characterGenerator[1881] = 8'hcc;
assign _c_characterGenerator[1882] = 8'hcc;
assign _c_characterGenerator[1883] = 8'h76;
assign _c_characterGenerator[1884] = 8'h00;
assign _c_characterGenerator[1885] = 8'h00;
assign _c_characterGenerator[1886] = 8'h00;
assign _c_characterGenerator[1887] = 8'h00;
assign _c_characterGenerator[1888] = 8'h00;
assign _c_characterGenerator[1889] = 8'h00;
assign _c_characterGenerator[1890] = 8'h00;
assign _c_characterGenerator[1891] = 8'h00;
assign _c_characterGenerator[1892] = 8'h00;
assign _c_characterGenerator[1893] = 8'h66;
assign _c_characterGenerator[1894] = 8'h66;
assign _c_characterGenerator[1895] = 8'h66;
assign _c_characterGenerator[1896] = 8'h66;
assign _c_characterGenerator[1897] = 8'h66;
assign _c_characterGenerator[1898] = 8'h3c;
assign _c_characterGenerator[1899] = 8'h18;
assign _c_characterGenerator[1900] = 8'h00;
assign _c_characterGenerator[1901] = 8'h00;
assign _c_characterGenerator[1902] = 8'h00;
assign _c_characterGenerator[1903] = 8'h00;
assign _c_characterGenerator[1904] = 8'h00;
assign _c_characterGenerator[1905] = 8'h00;
assign _c_characterGenerator[1906] = 8'h00;
assign _c_characterGenerator[1907] = 8'h00;
assign _c_characterGenerator[1908] = 8'h00;
assign _c_characterGenerator[1909] = 8'hc6;
assign _c_characterGenerator[1910] = 8'hc6;
assign _c_characterGenerator[1911] = 8'hd6;
assign _c_characterGenerator[1912] = 8'hd6;
assign _c_characterGenerator[1913] = 8'hd6;
assign _c_characterGenerator[1914] = 8'hfe;
assign _c_characterGenerator[1915] = 8'h6c;
assign _c_characterGenerator[1916] = 8'h00;
assign _c_characterGenerator[1917] = 8'h00;
assign _c_characterGenerator[1918] = 8'h00;
assign _c_characterGenerator[1919] = 8'h00;
assign _c_characterGenerator[1920] = 8'h00;
assign _c_characterGenerator[1921] = 8'h00;
assign _c_characterGenerator[1922] = 8'h00;
assign _c_characterGenerator[1923] = 8'h00;
assign _c_characterGenerator[1924] = 8'h00;
assign _c_characterGenerator[1925] = 8'hc6;
assign _c_characterGenerator[1926] = 8'h6c;
assign _c_characterGenerator[1927] = 8'h38;
assign _c_characterGenerator[1928] = 8'h38;
assign _c_characterGenerator[1929] = 8'h38;
assign _c_characterGenerator[1930] = 8'h6c;
assign _c_characterGenerator[1931] = 8'hc6;
assign _c_characterGenerator[1932] = 8'h00;
assign _c_characterGenerator[1933] = 8'h00;
assign _c_characterGenerator[1934] = 8'h00;
assign _c_characterGenerator[1935] = 8'h00;
assign _c_characterGenerator[1936] = 8'h00;
assign _c_characterGenerator[1937] = 8'h00;
assign _c_characterGenerator[1938] = 8'h00;
assign _c_characterGenerator[1939] = 8'h00;
assign _c_characterGenerator[1940] = 8'h00;
assign _c_characterGenerator[1941] = 8'hc6;
assign _c_characterGenerator[1942] = 8'hc6;
assign _c_characterGenerator[1943] = 8'hc6;
assign _c_characterGenerator[1944] = 8'hc6;
assign _c_characterGenerator[1945] = 8'hc6;
assign _c_characterGenerator[1946] = 8'hc6;
assign _c_characterGenerator[1947] = 8'h7e;
assign _c_characterGenerator[1948] = 8'h06;
assign _c_characterGenerator[1949] = 8'h0c;
assign _c_characterGenerator[1950] = 8'hf8;
assign _c_characterGenerator[1951] = 8'h00;
assign _c_characterGenerator[1952] = 8'h00;
assign _c_characterGenerator[1953] = 8'h00;
assign _c_characterGenerator[1954] = 8'h00;
assign _c_characterGenerator[1955] = 8'h00;
assign _c_characterGenerator[1956] = 8'h00;
assign _c_characterGenerator[1957] = 8'hfe;
assign _c_characterGenerator[1958] = 8'hcc;
assign _c_characterGenerator[1959] = 8'h18;
assign _c_characterGenerator[1960] = 8'h30;
assign _c_characterGenerator[1961] = 8'h60;
assign _c_characterGenerator[1962] = 8'hc6;
assign _c_characterGenerator[1963] = 8'hfe;
assign _c_characterGenerator[1964] = 8'h00;
assign _c_characterGenerator[1965] = 8'h00;
assign _c_characterGenerator[1966] = 8'h00;
assign _c_characterGenerator[1967] = 8'h00;
assign _c_characterGenerator[1968] = 8'h00;
assign _c_characterGenerator[1969] = 8'h00;
assign _c_characterGenerator[1970] = 8'h0e;
assign _c_characterGenerator[1971] = 8'h18;
assign _c_characterGenerator[1972] = 8'h18;
assign _c_characterGenerator[1973] = 8'h18;
assign _c_characterGenerator[1974] = 8'h70;
assign _c_characterGenerator[1975] = 8'h18;
assign _c_characterGenerator[1976] = 8'h18;
assign _c_characterGenerator[1977] = 8'h18;
assign _c_characterGenerator[1978] = 8'h18;
assign _c_characterGenerator[1979] = 8'h0e;
assign _c_characterGenerator[1980] = 8'h00;
assign _c_characterGenerator[1981] = 8'h00;
assign _c_characterGenerator[1982] = 8'h00;
assign _c_characterGenerator[1983] = 8'h00;
assign _c_characterGenerator[1984] = 8'h00;
assign _c_characterGenerator[1985] = 8'h00;
assign _c_characterGenerator[1986] = 8'h18;
assign _c_characterGenerator[1987] = 8'h18;
assign _c_characterGenerator[1988] = 8'h18;
assign _c_characterGenerator[1989] = 8'h18;
assign _c_characterGenerator[1990] = 8'h00;
assign _c_characterGenerator[1991] = 8'h18;
assign _c_characterGenerator[1992] = 8'h18;
assign _c_characterGenerator[1993] = 8'h18;
assign _c_characterGenerator[1994] = 8'h18;
assign _c_characterGenerator[1995] = 8'h18;
assign _c_characterGenerator[1996] = 8'h00;
assign _c_characterGenerator[1997] = 8'h00;
assign _c_characterGenerator[1998] = 8'h00;
assign _c_characterGenerator[1999] = 8'h00;
assign _c_characterGenerator[2000] = 8'h00;
assign _c_characterGenerator[2001] = 8'h00;
assign _c_characterGenerator[2002] = 8'h70;
assign _c_characterGenerator[2003] = 8'h18;
assign _c_characterGenerator[2004] = 8'h18;
assign _c_characterGenerator[2005] = 8'h18;
assign _c_characterGenerator[2006] = 8'h0e;
assign _c_characterGenerator[2007] = 8'h18;
assign _c_characterGenerator[2008] = 8'h18;
assign _c_characterGenerator[2009] = 8'h18;
assign _c_characterGenerator[2010] = 8'h18;
assign _c_characterGenerator[2011] = 8'h70;
assign _c_characterGenerator[2012] = 8'h00;
assign _c_characterGenerator[2013] = 8'h00;
assign _c_characterGenerator[2014] = 8'h00;
assign _c_characterGenerator[2015] = 8'h00;
assign _c_characterGenerator[2016] = 8'h00;
assign _c_characterGenerator[2017] = 8'h00;
assign _c_characterGenerator[2018] = 8'h76;
assign _c_characterGenerator[2019] = 8'hdc;
assign _c_characterGenerator[2020] = 8'h00;
assign _c_characterGenerator[2021] = 8'h00;
assign _c_characterGenerator[2022] = 8'h00;
assign _c_characterGenerator[2023] = 8'h00;
assign _c_characterGenerator[2024] = 8'h00;
assign _c_characterGenerator[2025] = 8'h00;
assign _c_characterGenerator[2026] = 8'h00;
assign _c_characterGenerator[2027] = 8'h00;
assign _c_characterGenerator[2028] = 8'h00;
assign _c_characterGenerator[2029] = 8'h00;
assign _c_characterGenerator[2030] = 8'h00;
assign _c_characterGenerator[2031] = 8'h00;
assign _c_characterGenerator[2032] = 8'h00;
assign _c_characterGenerator[2033] = 8'h00;
assign _c_characterGenerator[2034] = 8'h00;
assign _c_characterGenerator[2035] = 8'h00;
assign _c_characterGenerator[2036] = 8'h10;
assign _c_characterGenerator[2037] = 8'h38;
assign _c_characterGenerator[2038] = 8'h6c;
assign _c_characterGenerator[2039] = 8'hc6;
assign _c_characterGenerator[2040] = 8'hc6;
assign _c_characterGenerator[2041] = 8'hc6;
assign _c_characterGenerator[2042] = 8'hfe;
assign _c_characterGenerator[2043] = 8'h00;
assign _c_characterGenerator[2044] = 8'h00;
assign _c_characterGenerator[2045] = 8'h00;
assign _c_characterGenerator[2046] = 8'h00;
assign _c_characterGenerator[2047] = 8'h00;
assign _c_characterGenerator[2048] = 8'h00;
assign _c_characterGenerator[2049] = 8'h00;
assign _c_characterGenerator[2050] = 8'h3c;
assign _c_characterGenerator[2051] = 8'h66;
assign _c_characterGenerator[2052] = 8'hc2;
assign _c_characterGenerator[2053] = 8'hc0;
assign _c_characterGenerator[2054] = 8'hc0;
assign _c_characterGenerator[2055] = 8'hc0;
assign _c_characterGenerator[2056] = 8'hc2;
assign _c_characterGenerator[2057] = 8'h66;
assign _c_characterGenerator[2058] = 8'h3c;
assign _c_characterGenerator[2059] = 8'h0c;
assign _c_characterGenerator[2060] = 8'h06;
assign _c_characterGenerator[2061] = 8'h7c;
assign _c_characterGenerator[2062] = 8'h00;
assign _c_characterGenerator[2063] = 8'h00;
assign _c_characterGenerator[2064] = 8'h00;
assign _c_characterGenerator[2065] = 8'h00;
assign _c_characterGenerator[2066] = 8'hcc;
assign _c_characterGenerator[2067] = 8'h00;
assign _c_characterGenerator[2068] = 8'h00;
assign _c_characterGenerator[2069] = 8'hcc;
assign _c_characterGenerator[2070] = 8'hcc;
assign _c_characterGenerator[2071] = 8'hcc;
assign _c_characterGenerator[2072] = 8'hcc;
assign _c_characterGenerator[2073] = 8'hcc;
assign _c_characterGenerator[2074] = 8'hcc;
assign _c_characterGenerator[2075] = 8'h76;
assign _c_characterGenerator[2076] = 8'h00;
assign _c_characterGenerator[2077] = 8'h00;
assign _c_characterGenerator[2078] = 8'h00;
assign _c_characterGenerator[2079] = 8'h00;
assign _c_characterGenerator[2080] = 8'h00;
assign _c_characterGenerator[2081] = 8'h0c;
assign _c_characterGenerator[2082] = 8'h18;
assign _c_characterGenerator[2083] = 8'h30;
assign _c_characterGenerator[2084] = 8'h00;
assign _c_characterGenerator[2085] = 8'h7c;
assign _c_characterGenerator[2086] = 8'hc6;
assign _c_characterGenerator[2087] = 8'hfe;
assign _c_characterGenerator[2088] = 8'hc0;
assign _c_characterGenerator[2089] = 8'hc0;
assign _c_characterGenerator[2090] = 8'hc6;
assign _c_characterGenerator[2091] = 8'h7c;
assign _c_characterGenerator[2092] = 8'h00;
assign _c_characterGenerator[2093] = 8'h00;
assign _c_characterGenerator[2094] = 8'h00;
assign _c_characterGenerator[2095] = 8'h00;
assign _c_characterGenerator[2096] = 8'h00;
assign _c_characterGenerator[2097] = 8'h10;
assign _c_characterGenerator[2098] = 8'h38;
assign _c_characterGenerator[2099] = 8'h6c;
assign _c_characterGenerator[2100] = 8'h00;
assign _c_characterGenerator[2101] = 8'h78;
assign _c_characterGenerator[2102] = 8'h0c;
assign _c_characterGenerator[2103] = 8'h7c;
assign _c_characterGenerator[2104] = 8'hcc;
assign _c_characterGenerator[2105] = 8'hcc;
assign _c_characterGenerator[2106] = 8'hcc;
assign _c_characterGenerator[2107] = 8'h76;
assign _c_characterGenerator[2108] = 8'h00;
assign _c_characterGenerator[2109] = 8'h00;
assign _c_characterGenerator[2110] = 8'h00;
assign _c_characterGenerator[2111] = 8'h00;
assign _c_characterGenerator[2112] = 8'h00;
assign _c_characterGenerator[2113] = 8'h00;
assign _c_characterGenerator[2114] = 8'hcc;
assign _c_characterGenerator[2115] = 8'h00;
assign _c_characterGenerator[2116] = 8'h00;
assign _c_characterGenerator[2117] = 8'h78;
assign _c_characterGenerator[2118] = 8'h0c;
assign _c_characterGenerator[2119] = 8'h7c;
assign _c_characterGenerator[2120] = 8'hcc;
assign _c_characterGenerator[2121] = 8'hcc;
assign _c_characterGenerator[2122] = 8'hcc;
assign _c_characterGenerator[2123] = 8'h76;
assign _c_characterGenerator[2124] = 8'h00;
assign _c_characterGenerator[2125] = 8'h00;
assign _c_characterGenerator[2126] = 8'h00;
assign _c_characterGenerator[2127] = 8'h00;
assign _c_characterGenerator[2128] = 8'h00;
assign _c_characterGenerator[2129] = 8'h60;
assign _c_characterGenerator[2130] = 8'h30;
assign _c_characterGenerator[2131] = 8'h18;
assign _c_characterGenerator[2132] = 8'h00;
assign _c_characterGenerator[2133] = 8'h78;
assign _c_characterGenerator[2134] = 8'h0c;
assign _c_characterGenerator[2135] = 8'h7c;
assign _c_characterGenerator[2136] = 8'hcc;
assign _c_characterGenerator[2137] = 8'hcc;
assign _c_characterGenerator[2138] = 8'hcc;
assign _c_characterGenerator[2139] = 8'h76;
assign _c_characterGenerator[2140] = 8'h00;
assign _c_characterGenerator[2141] = 8'h00;
assign _c_characterGenerator[2142] = 8'h00;
assign _c_characterGenerator[2143] = 8'h00;
assign _c_characterGenerator[2144] = 8'h00;
assign _c_characterGenerator[2145] = 8'h38;
assign _c_characterGenerator[2146] = 8'h6c;
assign _c_characterGenerator[2147] = 8'h38;
assign _c_characterGenerator[2148] = 8'h00;
assign _c_characterGenerator[2149] = 8'h78;
assign _c_characterGenerator[2150] = 8'h0c;
assign _c_characterGenerator[2151] = 8'h7c;
assign _c_characterGenerator[2152] = 8'hcc;
assign _c_characterGenerator[2153] = 8'hcc;
assign _c_characterGenerator[2154] = 8'hcc;
assign _c_characterGenerator[2155] = 8'h76;
assign _c_characterGenerator[2156] = 8'h00;
assign _c_characterGenerator[2157] = 8'h00;
assign _c_characterGenerator[2158] = 8'h00;
assign _c_characterGenerator[2159] = 8'h00;
assign _c_characterGenerator[2160] = 8'h00;
assign _c_characterGenerator[2161] = 8'h00;
assign _c_characterGenerator[2162] = 8'h00;
assign _c_characterGenerator[2163] = 8'h00;
assign _c_characterGenerator[2164] = 8'h3c;
assign _c_characterGenerator[2165] = 8'h66;
assign _c_characterGenerator[2166] = 8'h60;
assign _c_characterGenerator[2167] = 8'h60;
assign _c_characterGenerator[2168] = 8'h66;
assign _c_characterGenerator[2169] = 8'h3c;
assign _c_characterGenerator[2170] = 8'h0c;
assign _c_characterGenerator[2171] = 8'h06;
assign _c_characterGenerator[2172] = 8'h3c;
assign _c_characterGenerator[2173] = 8'h00;
assign _c_characterGenerator[2174] = 8'h00;
assign _c_characterGenerator[2175] = 8'h00;
assign _c_characterGenerator[2176] = 8'h00;
assign _c_characterGenerator[2177] = 8'h10;
assign _c_characterGenerator[2178] = 8'h38;
assign _c_characterGenerator[2179] = 8'h6c;
assign _c_characterGenerator[2180] = 8'h00;
assign _c_characterGenerator[2181] = 8'h7c;
assign _c_characterGenerator[2182] = 8'hc6;
assign _c_characterGenerator[2183] = 8'hfe;
assign _c_characterGenerator[2184] = 8'hc0;
assign _c_characterGenerator[2185] = 8'hc0;
assign _c_characterGenerator[2186] = 8'hc6;
assign _c_characterGenerator[2187] = 8'h7c;
assign _c_characterGenerator[2188] = 8'h00;
assign _c_characterGenerator[2189] = 8'h00;
assign _c_characterGenerator[2190] = 8'h00;
assign _c_characterGenerator[2191] = 8'h00;
assign _c_characterGenerator[2192] = 8'h00;
assign _c_characterGenerator[2193] = 8'h00;
assign _c_characterGenerator[2194] = 8'hc6;
assign _c_characterGenerator[2195] = 8'h00;
assign _c_characterGenerator[2196] = 8'h00;
assign _c_characterGenerator[2197] = 8'h7c;
assign _c_characterGenerator[2198] = 8'hc6;
assign _c_characterGenerator[2199] = 8'hfe;
assign _c_characterGenerator[2200] = 8'hc0;
assign _c_characterGenerator[2201] = 8'hc0;
assign _c_characterGenerator[2202] = 8'hc6;
assign _c_characterGenerator[2203] = 8'h7c;
assign _c_characterGenerator[2204] = 8'h00;
assign _c_characterGenerator[2205] = 8'h00;
assign _c_characterGenerator[2206] = 8'h00;
assign _c_characterGenerator[2207] = 8'h00;
assign _c_characterGenerator[2208] = 8'h00;
assign _c_characterGenerator[2209] = 8'h60;
assign _c_characterGenerator[2210] = 8'h30;
assign _c_characterGenerator[2211] = 8'h18;
assign _c_characterGenerator[2212] = 8'h00;
assign _c_characterGenerator[2213] = 8'h7c;
assign _c_characterGenerator[2214] = 8'hc6;
assign _c_characterGenerator[2215] = 8'hfe;
assign _c_characterGenerator[2216] = 8'hc0;
assign _c_characterGenerator[2217] = 8'hc0;
assign _c_characterGenerator[2218] = 8'hc6;
assign _c_characterGenerator[2219] = 8'h7c;
assign _c_characterGenerator[2220] = 8'h00;
assign _c_characterGenerator[2221] = 8'h00;
assign _c_characterGenerator[2222] = 8'h00;
assign _c_characterGenerator[2223] = 8'h00;
assign _c_characterGenerator[2224] = 8'h00;
assign _c_characterGenerator[2225] = 8'h00;
assign _c_characterGenerator[2226] = 8'h66;
assign _c_characterGenerator[2227] = 8'h00;
assign _c_characterGenerator[2228] = 8'h00;
assign _c_characterGenerator[2229] = 8'h38;
assign _c_characterGenerator[2230] = 8'h18;
assign _c_characterGenerator[2231] = 8'h18;
assign _c_characterGenerator[2232] = 8'h18;
assign _c_characterGenerator[2233] = 8'h18;
assign _c_characterGenerator[2234] = 8'h18;
assign _c_characterGenerator[2235] = 8'h3c;
assign _c_characterGenerator[2236] = 8'h00;
assign _c_characterGenerator[2237] = 8'h00;
assign _c_characterGenerator[2238] = 8'h00;
assign _c_characterGenerator[2239] = 8'h00;
assign _c_characterGenerator[2240] = 8'h00;
assign _c_characterGenerator[2241] = 8'h18;
assign _c_characterGenerator[2242] = 8'h3c;
assign _c_characterGenerator[2243] = 8'h66;
assign _c_characterGenerator[2244] = 8'h00;
assign _c_characterGenerator[2245] = 8'h38;
assign _c_characterGenerator[2246] = 8'h18;
assign _c_characterGenerator[2247] = 8'h18;
assign _c_characterGenerator[2248] = 8'h18;
assign _c_characterGenerator[2249] = 8'h18;
assign _c_characterGenerator[2250] = 8'h18;
assign _c_characterGenerator[2251] = 8'h3c;
assign _c_characterGenerator[2252] = 8'h00;
assign _c_characterGenerator[2253] = 8'h00;
assign _c_characterGenerator[2254] = 8'h00;
assign _c_characterGenerator[2255] = 8'h00;
assign _c_characterGenerator[2256] = 8'h00;
assign _c_characterGenerator[2257] = 8'h60;
assign _c_characterGenerator[2258] = 8'h30;
assign _c_characterGenerator[2259] = 8'h18;
assign _c_characterGenerator[2260] = 8'h00;
assign _c_characterGenerator[2261] = 8'h38;
assign _c_characterGenerator[2262] = 8'h18;
assign _c_characterGenerator[2263] = 8'h18;
assign _c_characterGenerator[2264] = 8'h18;
assign _c_characterGenerator[2265] = 8'h18;
assign _c_characterGenerator[2266] = 8'h18;
assign _c_characterGenerator[2267] = 8'h3c;
assign _c_characterGenerator[2268] = 8'h00;
assign _c_characterGenerator[2269] = 8'h00;
assign _c_characterGenerator[2270] = 8'h00;
assign _c_characterGenerator[2271] = 8'h00;
assign _c_characterGenerator[2272] = 8'h00;
assign _c_characterGenerator[2273] = 8'hc6;
assign _c_characterGenerator[2274] = 8'h00;
assign _c_characterGenerator[2275] = 8'h10;
assign _c_characterGenerator[2276] = 8'h38;
assign _c_characterGenerator[2277] = 8'h6c;
assign _c_characterGenerator[2278] = 8'hc6;
assign _c_characterGenerator[2279] = 8'hc6;
assign _c_characterGenerator[2280] = 8'hfe;
assign _c_characterGenerator[2281] = 8'hc6;
assign _c_characterGenerator[2282] = 8'hc6;
assign _c_characterGenerator[2283] = 8'hc6;
assign _c_characterGenerator[2284] = 8'h00;
assign _c_characterGenerator[2285] = 8'h00;
assign _c_characterGenerator[2286] = 8'h00;
assign _c_characterGenerator[2287] = 8'h00;
assign _c_characterGenerator[2288] = 8'h38;
assign _c_characterGenerator[2289] = 8'h6c;
assign _c_characterGenerator[2290] = 8'h38;
assign _c_characterGenerator[2291] = 8'h00;
assign _c_characterGenerator[2292] = 8'h38;
assign _c_characterGenerator[2293] = 8'h6c;
assign _c_characterGenerator[2294] = 8'hc6;
assign _c_characterGenerator[2295] = 8'hc6;
assign _c_characterGenerator[2296] = 8'hfe;
assign _c_characterGenerator[2297] = 8'hc6;
assign _c_characterGenerator[2298] = 8'hc6;
assign _c_characterGenerator[2299] = 8'hc6;
assign _c_characterGenerator[2300] = 8'h00;
assign _c_characterGenerator[2301] = 8'h00;
assign _c_characterGenerator[2302] = 8'h00;
assign _c_characterGenerator[2303] = 8'h00;
assign _c_characterGenerator[2304] = 8'h18;
assign _c_characterGenerator[2305] = 8'h30;
assign _c_characterGenerator[2306] = 8'h60;
assign _c_characterGenerator[2307] = 8'h00;
assign _c_characterGenerator[2308] = 8'hfe;
assign _c_characterGenerator[2309] = 8'h66;
assign _c_characterGenerator[2310] = 8'h60;
assign _c_characterGenerator[2311] = 8'h7c;
assign _c_characterGenerator[2312] = 8'h60;
assign _c_characterGenerator[2313] = 8'h60;
assign _c_characterGenerator[2314] = 8'h66;
assign _c_characterGenerator[2315] = 8'hfe;
assign _c_characterGenerator[2316] = 8'h00;
assign _c_characterGenerator[2317] = 8'h00;
assign _c_characterGenerator[2318] = 8'h00;
assign _c_characterGenerator[2319] = 8'h00;
assign _c_characterGenerator[2320] = 8'h00;
assign _c_characterGenerator[2321] = 8'h00;
assign _c_characterGenerator[2322] = 8'h00;
assign _c_characterGenerator[2323] = 8'h00;
assign _c_characterGenerator[2324] = 8'h00;
assign _c_characterGenerator[2325] = 8'hcc;
assign _c_characterGenerator[2326] = 8'h76;
assign _c_characterGenerator[2327] = 8'h36;
assign _c_characterGenerator[2328] = 8'h7e;
assign _c_characterGenerator[2329] = 8'hd8;
assign _c_characterGenerator[2330] = 8'hd8;
assign _c_characterGenerator[2331] = 8'h6e;
assign _c_characterGenerator[2332] = 8'h00;
assign _c_characterGenerator[2333] = 8'h00;
assign _c_characterGenerator[2334] = 8'h00;
assign _c_characterGenerator[2335] = 8'h00;
assign _c_characterGenerator[2336] = 8'h00;
assign _c_characterGenerator[2337] = 8'h00;
assign _c_characterGenerator[2338] = 8'h3e;
assign _c_characterGenerator[2339] = 8'h6c;
assign _c_characterGenerator[2340] = 8'hcc;
assign _c_characterGenerator[2341] = 8'hcc;
assign _c_characterGenerator[2342] = 8'hfe;
assign _c_characterGenerator[2343] = 8'hcc;
assign _c_characterGenerator[2344] = 8'hcc;
assign _c_characterGenerator[2345] = 8'hcc;
assign _c_characterGenerator[2346] = 8'hcc;
assign _c_characterGenerator[2347] = 8'hce;
assign _c_characterGenerator[2348] = 8'h00;
assign _c_characterGenerator[2349] = 8'h00;
assign _c_characterGenerator[2350] = 8'h00;
assign _c_characterGenerator[2351] = 8'h00;
assign _c_characterGenerator[2352] = 8'h00;
assign _c_characterGenerator[2353] = 8'h10;
assign _c_characterGenerator[2354] = 8'h38;
assign _c_characterGenerator[2355] = 8'h6c;
assign _c_characterGenerator[2356] = 8'h00;
assign _c_characterGenerator[2357] = 8'h7c;
assign _c_characterGenerator[2358] = 8'hc6;
assign _c_characterGenerator[2359] = 8'hc6;
assign _c_characterGenerator[2360] = 8'hc6;
assign _c_characterGenerator[2361] = 8'hc6;
assign _c_characterGenerator[2362] = 8'hc6;
assign _c_characterGenerator[2363] = 8'h7c;
assign _c_characterGenerator[2364] = 8'h00;
assign _c_characterGenerator[2365] = 8'h00;
assign _c_characterGenerator[2366] = 8'h00;
assign _c_characterGenerator[2367] = 8'h00;
assign _c_characterGenerator[2368] = 8'h00;
assign _c_characterGenerator[2369] = 8'h00;
assign _c_characterGenerator[2370] = 8'hc6;
assign _c_characterGenerator[2371] = 8'h00;
assign _c_characterGenerator[2372] = 8'h00;
assign _c_characterGenerator[2373] = 8'h7c;
assign _c_characterGenerator[2374] = 8'hc6;
assign _c_characterGenerator[2375] = 8'hc6;
assign _c_characterGenerator[2376] = 8'hc6;
assign _c_characterGenerator[2377] = 8'hc6;
assign _c_characterGenerator[2378] = 8'hc6;
assign _c_characterGenerator[2379] = 8'h7c;
assign _c_characterGenerator[2380] = 8'h00;
assign _c_characterGenerator[2381] = 8'h00;
assign _c_characterGenerator[2382] = 8'h00;
assign _c_characterGenerator[2383] = 8'h00;
assign _c_characterGenerator[2384] = 8'h00;
assign _c_characterGenerator[2385] = 8'h60;
assign _c_characterGenerator[2386] = 8'h30;
assign _c_characterGenerator[2387] = 8'h18;
assign _c_characterGenerator[2388] = 8'h00;
assign _c_characterGenerator[2389] = 8'h7c;
assign _c_characterGenerator[2390] = 8'hc6;
assign _c_characterGenerator[2391] = 8'hc6;
assign _c_characterGenerator[2392] = 8'hc6;
assign _c_characterGenerator[2393] = 8'hc6;
assign _c_characterGenerator[2394] = 8'hc6;
assign _c_characterGenerator[2395] = 8'h7c;
assign _c_characterGenerator[2396] = 8'h00;
assign _c_characterGenerator[2397] = 8'h00;
assign _c_characterGenerator[2398] = 8'h00;
assign _c_characterGenerator[2399] = 8'h00;
assign _c_characterGenerator[2400] = 8'h00;
assign _c_characterGenerator[2401] = 8'h30;
assign _c_characterGenerator[2402] = 8'h78;
assign _c_characterGenerator[2403] = 8'hcc;
assign _c_characterGenerator[2404] = 8'h00;
assign _c_characterGenerator[2405] = 8'hcc;
assign _c_characterGenerator[2406] = 8'hcc;
assign _c_characterGenerator[2407] = 8'hcc;
assign _c_characterGenerator[2408] = 8'hcc;
assign _c_characterGenerator[2409] = 8'hcc;
assign _c_characterGenerator[2410] = 8'hcc;
assign _c_characterGenerator[2411] = 8'h76;
assign _c_characterGenerator[2412] = 8'h00;
assign _c_characterGenerator[2413] = 8'h00;
assign _c_characterGenerator[2414] = 8'h00;
assign _c_characterGenerator[2415] = 8'h00;
assign _c_characterGenerator[2416] = 8'h00;
assign _c_characterGenerator[2417] = 8'h60;
assign _c_characterGenerator[2418] = 8'h30;
assign _c_characterGenerator[2419] = 8'h18;
assign _c_characterGenerator[2420] = 8'h00;
assign _c_characterGenerator[2421] = 8'hcc;
assign _c_characterGenerator[2422] = 8'hcc;
assign _c_characterGenerator[2423] = 8'hcc;
assign _c_characterGenerator[2424] = 8'hcc;
assign _c_characterGenerator[2425] = 8'hcc;
assign _c_characterGenerator[2426] = 8'hcc;
assign _c_characterGenerator[2427] = 8'h76;
assign _c_characterGenerator[2428] = 8'h00;
assign _c_characterGenerator[2429] = 8'h00;
assign _c_characterGenerator[2430] = 8'h00;
assign _c_characterGenerator[2431] = 8'h00;
assign _c_characterGenerator[2432] = 8'h00;
assign _c_characterGenerator[2433] = 8'h00;
assign _c_characterGenerator[2434] = 8'hc6;
assign _c_characterGenerator[2435] = 8'h00;
assign _c_characterGenerator[2436] = 8'h00;
assign _c_characterGenerator[2437] = 8'hc6;
assign _c_characterGenerator[2438] = 8'hc6;
assign _c_characterGenerator[2439] = 8'hc6;
assign _c_characterGenerator[2440] = 8'hc6;
assign _c_characterGenerator[2441] = 8'hc6;
assign _c_characterGenerator[2442] = 8'hc6;
assign _c_characterGenerator[2443] = 8'h7e;
assign _c_characterGenerator[2444] = 8'h06;
assign _c_characterGenerator[2445] = 8'h0c;
assign _c_characterGenerator[2446] = 8'h78;
assign _c_characterGenerator[2447] = 8'h00;
assign _c_characterGenerator[2448] = 8'h00;
assign _c_characterGenerator[2449] = 8'hc6;
assign _c_characterGenerator[2450] = 8'h00;
assign _c_characterGenerator[2451] = 8'h7c;
assign _c_characterGenerator[2452] = 8'hc6;
assign _c_characterGenerator[2453] = 8'hc6;
assign _c_characterGenerator[2454] = 8'hc6;
assign _c_characterGenerator[2455] = 8'hc6;
assign _c_characterGenerator[2456] = 8'hc6;
assign _c_characterGenerator[2457] = 8'hc6;
assign _c_characterGenerator[2458] = 8'hc6;
assign _c_characterGenerator[2459] = 8'h7c;
assign _c_characterGenerator[2460] = 8'h00;
assign _c_characterGenerator[2461] = 8'h00;
assign _c_characterGenerator[2462] = 8'h00;
assign _c_characterGenerator[2463] = 8'h00;
assign _c_characterGenerator[2464] = 8'h00;
assign _c_characterGenerator[2465] = 8'hc6;
assign _c_characterGenerator[2466] = 8'h00;
assign _c_characterGenerator[2467] = 8'hc6;
assign _c_characterGenerator[2468] = 8'hc6;
assign _c_characterGenerator[2469] = 8'hc6;
assign _c_characterGenerator[2470] = 8'hc6;
assign _c_characterGenerator[2471] = 8'hc6;
assign _c_characterGenerator[2472] = 8'hc6;
assign _c_characterGenerator[2473] = 8'hc6;
assign _c_characterGenerator[2474] = 8'hc6;
assign _c_characterGenerator[2475] = 8'h7c;
assign _c_characterGenerator[2476] = 8'h00;
assign _c_characterGenerator[2477] = 8'h00;
assign _c_characterGenerator[2478] = 8'h00;
assign _c_characterGenerator[2479] = 8'h00;
assign _c_characterGenerator[2480] = 8'h00;
assign _c_characterGenerator[2481] = 8'h18;
assign _c_characterGenerator[2482] = 8'h18;
assign _c_characterGenerator[2483] = 8'h3c;
assign _c_characterGenerator[2484] = 8'h66;
assign _c_characterGenerator[2485] = 8'h60;
assign _c_characterGenerator[2486] = 8'h60;
assign _c_characterGenerator[2487] = 8'h60;
assign _c_characterGenerator[2488] = 8'h66;
assign _c_characterGenerator[2489] = 8'h3c;
assign _c_characterGenerator[2490] = 8'h18;
assign _c_characterGenerator[2491] = 8'h18;
assign _c_characterGenerator[2492] = 8'h00;
assign _c_characterGenerator[2493] = 8'h00;
assign _c_characterGenerator[2494] = 8'h00;
assign _c_characterGenerator[2495] = 8'h00;
assign _c_characterGenerator[2496] = 8'h00;
assign _c_characterGenerator[2497] = 8'h38;
assign _c_characterGenerator[2498] = 8'h6c;
assign _c_characterGenerator[2499] = 8'h64;
assign _c_characterGenerator[2500] = 8'h60;
assign _c_characterGenerator[2501] = 8'hf0;
assign _c_characterGenerator[2502] = 8'h60;
assign _c_characterGenerator[2503] = 8'h60;
assign _c_characterGenerator[2504] = 8'h60;
assign _c_characterGenerator[2505] = 8'h60;
assign _c_characterGenerator[2506] = 8'he6;
assign _c_characterGenerator[2507] = 8'hfc;
assign _c_characterGenerator[2508] = 8'h00;
assign _c_characterGenerator[2509] = 8'h00;
assign _c_characterGenerator[2510] = 8'h00;
assign _c_characterGenerator[2511] = 8'h00;
assign _c_characterGenerator[2512] = 8'h00;
assign _c_characterGenerator[2513] = 8'h00;
assign _c_characterGenerator[2514] = 8'h66;
assign _c_characterGenerator[2515] = 8'h66;
assign _c_characterGenerator[2516] = 8'h3c;
assign _c_characterGenerator[2517] = 8'h18;
assign _c_characterGenerator[2518] = 8'h7e;
assign _c_characterGenerator[2519] = 8'h18;
assign _c_characterGenerator[2520] = 8'h7e;
assign _c_characterGenerator[2521] = 8'h18;
assign _c_characterGenerator[2522] = 8'h18;
assign _c_characterGenerator[2523] = 8'h18;
assign _c_characterGenerator[2524] = 8'h00;
assign _c_characterGenerator[2525] = 8'h00;
assign _c_characterGenerator[2526] = 8'h00;
assign _c_characterGenerator[2527] = 8'h00;
assign _c_characterGenerator[2528] = 8'h00;
assign _c_characterGenerator[2529] = 8'hf8;
assign _c_characterGenerator[2530] = 8'hcc;
assign _c_characterGenerator[2531] = 8'hcc;
assign _c_characterGenerator[2532] = 8'hf8;
assign _c_characterGenerator[2533] = 8'hc4;
assign _c_characterGenerator[2534] = 8'hcc;
assign _c_characterGenerator[2535] = 8'hde;
assign _c_characterGenerator[2536] = 8'hcc;
assign _c_characterGenerator[2537] = 8'hcc;
assign _c_characterGenerator[2538] = 8'hcc;
assign _c_characterGenerator[2539] = 8'hc6;
assign _c_characterGenerator[2540] = 8'h00;
assign _c_characterGenerator[2541] = 8'h00;
assign _c_characterGenerator[2542] = 8'h00;
assign _c_characterGenerator[2543] = 8'h00;
assign _c_characterGenerator[2544] = 8'h00;
assign _c_characterGenerator[2545] = 8'h0e;
assign _c_characterGenerator[2546] = 8'h1b;
assign _c_characterGenerator[2547] = 8'h18;
assign _c_characterGenerator[2548] = 8'h18;
assign _c_characterGenerator[2549] = 8'h18;
assign _c_characterGenerator[2550] = 8'h7e;
assign _c_characterGenerator[2551] = 8'h18;
assign _c_characterGenerator[2552] = 8'h18;
assign _c_characterGenerator[2553] = 8'h18;
assign _c_characterGenerator[2554] = 8'h18;
assign _c_characterGenerator[2555] = 8'h18;
assign _c_characterGenerator[2556] = 8'hd8;
assign _c_characterGenerator[2557] = 8'h70;
assign _c_characterGenerator[2558] = 8'h00;
assign _c_characterGenerator[2559] = 8'h00;
assign _c_characterGenerator[2560] = 8'h00;
assign _c_characterGenerator[2561] = 8'h18;
assign _c_characterGenerator[2562] = 8'h30;
assign _c_characterGenerator[2563] = 8'h60;
assign _c_characterGenerator[2564] = 8'h00;
assign _c_characterGenerator[2565] = 8'h78;
assign _c_characterGenerator[2566] = 8'h0c;
assign _c_characterGenerator[2567] = 8'h7c;
assign _c_characterGenerator[2568] = 8'hcc;
assign _c_characterGenerator[2569] = 8'hcc;
assign _c_characterGenerator[2570] = 8'hcc;
assign _c_characterGenerator[2571] = 8'h76;
assign _c_characterGenerator[2572] = 8'h00;
assign _c_characterGenerator[2573] = 8'h00;
assign _c_characterGenerator[2574] = 8'h00;
assign _c_characterGenerator[2575] = 8'h00;
assign _c_characterGenerator[2576] = 8'h00;
assign _c_characterGenerator[2577] = 8'h0c;
assign _c_characterGenerator[2578] = 8'h18;
assign _c_characterGenerator[2579] = 8'h30;
assign _c_characterGenerator[2580] = 8'h00;
assign _c_characterGenerator[2581] = 8'h38;
assign _c_characterGenerator[2582] = 8'h18;
assign _c_characterGenerator[2583] = 8'h18;
assign _c_characterGenerator[2584] = 8'h18;
assign _c_characterGenerator[2585] = 8'h18;
assign _c_characterGenerator[2586] = 8'h18;
assign _c_characterGenerator[2587] = 8'h3c;
assign _c_characterGenerator[2588] = 8'h00;
assign _c_characterGenerator[2589] = 8'h00;
assign _c_characterGenerator[2590] = 8'h00;
assign _c_characterGenerator[2591] = 8'h00;
assign _c_characterGenerator[2592] = 8'h00;
assign _c_characterGenerator[2593] = 8'h18;
assign _c_characterGenerator[2594] = 8'h30;
assign _c_characterGenerator[2595] = 8'h60;
assign _c_characterGenerator[2596] = 8'h00;
assign _c_characterGenerator[2597] = 8'h7c;
assign _c_characterGenerator[2598] = 8'hc6;
assign _c_characterGenerator[2599] = 8'hc6;
assign _c_characterGenerator[2600] = 8'hc6;
assign _c_characterGenerator[2601] = 8'hc6;
assign _c_characterGenerator[2602] = 8'hc6;
assign _c_characterGenerator[2603] = 8'h7c;
assign _c_characterGenerator[2604] = 8'h00;
assign _c_characterGenerator[2605] = 8'h00;
assign _c_characterGenerator[2606] = 8'h00;
assign _c_characterGenerator[2607] = 8'h00;
assign _c_characterGenerator[2608] = 8'h00;
assign _c_characterGenerator[2609] = 8'h18;
assign _c_characterGenerator[2610] = 8'h30;
assign _c_characterGenerator[2611] = 8'h60;
assign _c_characterGenerator[2612] = 8'h00;
assign _c_characterGenerator[2613] = 8'hcc;
assign _c_characterGenerator[2614] = 8'hcc;
assign _c_characterGenerator[2615] = 8'hcc;
assign _c_characterGenerator[2616] = 8'hcc;
assign _c_characterGenerator[2617] = 8'hcc;
assign _c_characterGenerator[2618] = 8'hcc;
assign _c_characterGenerator[2619] = 8'h76;
assign _c_characterGenerator[2620] = 8'h00;
assign _c_characterGenerator[2621] = 8'h00;
assign _c_characterGenerator[2622] = 8'h00;
assign _c_characterGenerator[2623] = 8'h00;
assign _c_characterGenerator[2624] = 8'h00;
assign _c_characterGenerator[2625] = 8'h00;
assign _c_characterGenerator[2626] = 8'h76;
assign _c_characterGenerator[2627] = 8'hdc;
assign _c_characterGenerator[2628] = 8'h00;
assign _c_characterGenerator[2629] = 8'hdc;
assign _c_characterGenerator[2630] = 8'h66;
assign _c_characterGenerator[2631] = 8'h66;
assign _c_characterGenerator[2632] = 8'h66;
assign _c_characterGenerator[2633] = 8'h66;
assign _c_characterGenerator[2634] = 8'h66;
assign _c_characterGenerator[2635] = 8'h66;
assign _c_characterGenerator[2636] = 8'h00;
assign _c_characterGenerator[2637] = 8'h00;
assign _c_characterGenerator[2638] = 8'h00;
assign _c_characterGenerator[2639] = 8'h00;
assign _c_characterGenerator[2640] = 8'h76;
assign _c_characterGenerator[2641] = 8'hdc;
assign _c_characterGenerator[2642] = 8'h00;
assign _c_characterGenerator[2643] = 8'hc6;
assign _c_characterGenerator[2644] = 8'he6;
assign _c_characterGenerator[2645] = 8'hf6;
assign _c_characterGenerator[2646] = 8'hfe;
assign _c_characterGenerator[2647] = 8'hde;
assign _c_characterGenerator[2648] = 8'hce;
assign _c_characterGenerator[2649] = 8'hc6;
assign _c_characterGenerator[2650] = 8'hc6;
assign _c_characterGenerator[2651] = 8'hc6;
assign _c_characterGenerator[2652] = 8'h00;
assign _c_characterGenerator[2653] = 8'h00;
assign _c_characterGenerator[2654] = 8'h00;
assign _c_characterGenerator[2655] = 8'h00;
assign _c_characterGenerator[2656] = 8'h00;
assign _c_characterGenerator[2657] = 8'h3c;
assign _c_characterGenerator[2658] = 8'h6c;
assign _c_characterGenerator[2659] = 8'h6c;
assign _c_characterGenerator[2660] = 8'h3e;
assign _c_characterGenerator[2661] = 8'h00;
assign _c_characterGenerator[2662] = 8'h7e;
assign _c_characterGenerator[2663] = 8'h00;
assign _c_characterGenerator[2664] = 8'h00;
assign _c_characterGenerator[2665] = 8'h00;
assign _c_characterGenerator[2666] = 8'h00;
assign _c_characterGenerator[2667] = 8'h00;
assign _c_characterGenerator[2668] = 8'h00;
assign _c_characterGenerator[2669] = 8'h00;
assign _c_characterGenerator[2670] = 8'h00;
assign _c_characterGenerator[2671] = 8'h00;
assign _c_characterGenerator[2672] = 8'h00;
assign _c_characterGenerator[2673] = 8'h38;
assign _c_characterGenerator[2674] = 8'h6c;
assign _c_characterGenerator[2675] = 8'h6c;
assign _c_characterGenerator[2676] = 8'h38;
assign _c_characterGenerator[2677] = 8'h00;
assign _c_characterGenerator[2678] = 8'h7c;
assign _c_characterGenerator[2679] = 8'h00;
assign _c_characterGenerator[2680] = 8'h00;
assign _c_characterGenerator[2681] = 8'h00;
assign _c_characterGenerator[2682] = 8'h00;
assign _c_characterGenerator[2683] = 8'h00;
assign _c_characterGenerator[2684] = 8'h00;
assign _c_characterGenerator[2685] = 8'h00;
assign _c_characterGenerator[2686] = 8'h00;
assign _c_characterGenerator[2687] = 8'h00;
assign _c_characterGenerator[2688] = 8'h00;
assign _c_characterGenerator[2689] = 8'h00;
assign _c_characterGenerator[2690] = 8'h30;
assign _c_characterGenerator[2691] = 8'h30;
assign _c_characterGenerator[2692] = 8'h00;
assign _c_characterGenerator[2693] = 8'h30;
assign _c_characterGenerator[2694] = 8'h30;
assign _c_characterGenerator[2695] = 8'h60;
assign _c_characterGenerator[2696] = 8'hc0;
assign _c_characterGenerator[2697] = 8'hc6;
assign _c_characterGenerator[2698] = 8'hc6;
assign _c_characterGenerator[2699] = 8'h7c;
assign _c_characterGenerator[2700] = 8'h00;
assign _c_characterGenerator[2701] = 8'h00;
assign _c_characterGenerator[2702] = 8'h00;
assign _c_characterGenerator[2703] = 8'h00;
assign _c_characterGenerator[2704] = 8'h00;
assign _c_characterGenerator[2705] = 8'h00;
assign _c_characterGenerator[2706] = 8'h00;
assign _c_characterGenerator[2707] = 8'h00;
assign _c_characterGenerator[2708] = 8'h00;
assign _c_characterGenerator[2709] = 8'h00;
assign _c_characterGenerator[2710] = 8'hfe;
assign _c_characterGenerator[2711] = 8'hc0;
assign _c_characterGenerator[2712] = 8'hc0;
assign _c_characterGenerator[2713] = 8'hc0;
assign _c_characterGenerator[2714] = 8'hc0;
assign _c_characterGenerator[2715] = 8'h00;
assign _c_characterGenerator[2716] = 8'h00;
assign _c_characterGenerator[2717] = 8'h00;
assign _c_characterGenerator[2718] = 8'h00;
assign _c_characterGenerator[2719] = 8'h00;
assign _c_characterGenerator[2720] = 8'h00;
assign _c_characterGenerator[2721] = 8'h00;
assign _c_characterGenerator[2722] = 8'h00;
assign _c_characterGenerator[2723] = 8'h00;
assign _c_characterGenerator[2724] = 8'h00;
assign _c_characterGenerator[2725] = 8'h00;
assign _c_characterGenerator[2726] = 8'hfe;
assign _c_characterGenerator[2727] = 8'h06;
assign _c_characterGenerator[2728] = 8'h06;
assign _c_characterGenerator[2729] = 8'h06;
assign _c_characterGenerator[2730] = 8'h06;
assign _c_characterGenerator[2731] = 8'h00;
assign _c_characterGenerator[2732] = 8'h00;
assign _c_characterGenerator[2733] = 8'h00;
assign _c_characterGenerator[2734] = 8'h00;
assign _c_characterGenerator[2735] = 8'h00;
assign _c_characterGenerator[2736] = 8'h00;
assign _c_characterGenerator[2737] = 8'hc0;
assign _c_characterGenerator[2738] = 8'hc0;
assign _c_characterGenerator[2739] = 8'hc2;
assign _c_characterGenerator[2740] = 8'hc6;
assign _c_characterGenerator[2741] = 8'hcc;
assign _c_characterGenerator[2742] = 8'h18;
assign _c_characterGenerator[2743] = 8'h30;
assign _c_characterGenerator[2744] = 8'h60;
assign _c_characterGenerator[2745] = 8'hdc;
assign _c_characterGenerator[2746] = 8'h86;
assign _c_characterGenerator[2747] = 8'h0c;
assign _c_characterGenerator[2748] = 8'h18;
assign _c_characterGenerator[2749] = 8'h3e;
assign _c_characterGenerator[2750] = 8'h00;
assign _c_characterGenerator[2751] = 8'h00;
assign _c_characterGenerator[2752] = 8'h00;
assign _c_characterGenerator[2753] = 8'hc0;
assign _c_characterGenerator[2754] = 8'hc0;
assign _c_characterGenerator[2755] = 8'hc2;
assign _c_characterGenerator[2756] = 8'hc6;
assign _c_characterGenerator[2757] = 8'hcc;
assign _c_characterGenerator[2758] = 8'h18;
assign _c_characterGenerator[2759] = 8'h30;
assign _c_characterGenerator[2760] = 8'h66;
assign _c_characterGenerator[2761] = 8'hce;
assign _c_characterGenerator[2762] = 8'h9e;
assign _c_characterGenerator[2763] = 8'h3e;
assign _c_characterGenerator[2764] = 8'h06;
assign _c_characterGenerator[2765] = 8'h06;
assign _c_characterGenerator[2766] = 8'h00;
assign _c_characterGenerator[2767] = 8'h00;
assign _c_characterGenerator[2768] = 8'h00;
assign _c_characterGenerator[2769] = 8'h00;
assign _c_characterGenerator[2770] = 8'h18;
assign _c_characterGenerator[2771] = 8'h18;
assign _c_characterGenerator[2772] = 8'h00;
assign _c_characterGenerator[2773] = 8'h18;
assign _c_characterGenerator[2774] = 8'h18;
assign _c_characterGenerator[2775] = 8'h18;
assign _c_characterGenerator[2776] = 8'h3c;
assign _c_characterGenerator[2777] = 8'h3c;
assign _c_characterGenerator[2778] = 8'h3c;
assign _c_characterGenerator[2779] = 8'h18;
assign _c_characterGenerator[2780] = 8'h00;
assign _c_characterGenerator[2781] = 8'h00;
assign _c_characterGenerator[2782] = 8'h00;
assign _c_characterGenerator[2783] = 8'h00;
assign _c_characterGenerator[2784] = 8'h00;
assign _c_characterGenerator[2785] = 8'h00;
assign _c_characterGenerator[2786] = 8'h00;
assign _c_characterGenerator[2787] = 8'h00;
assign _c_characterGenerator[2788] = 8'h00;
assign _c_characterGenerator[2789] = 8'h36;
assign _c_characterGenerator[2790] = 8'h6c;
assign _c_characterGenerator[2791] = 8'hd8;
assign _c_characterGenerator[2792] = 8'h6c;
assign _c_characterGenerator[2793] = 8'h36;
assign _c_characterGenerator[2794] = 8'h00;
assign _c_characterGenerator[2795] = 8'h00;
assign _c_characterGenerator[2796] = 8'h00;
assign _c_characterGenerator[2797] = 8'h00;
assign _c_characterGenerator[2798] = 8'h00;
assign _c_characterGenerator[2799] = 8'h00;
assign _c_characterGenerator[2800] = 8'h00;
assign _c_characterGenerator[2801] = 8'h00;
assign _c_characterGenerator[2802] = 8'h00;
assign _c_characterGenerator[2803] = 8'h00;
assign _c_characterGenerator[2804] = 8'h00;
assign _c_characterGenerator[2805] = 8'hd8;
assign _c_characterGenerator[2806] = 8'h6c;
assign _c_characterGenerator[2807] = 8'h36;
assign _c_characterGenerator[2808] = 8'h6c;
assign _c_characterGenerator[2809] = 8'hd8;
assign _c_characterGenerator[2810] = 8'h00;
assign _c_characterGenerator[2811] = 8'h00;
assign _c_characterGenerator[2812] = 8'h00;
assign _c_characterGenerator[2813] = 8'h00;
assign _c_characterGenerator[2814] = 8'h00;
assign _c_characterGenerator[2815] = 8'h00;
assign _c_characterGenerator[2816] = 8'h11;
assign _c_characterGenerator[2817] = 8'h44;
assign _c_characterGenerator[2818] = 8'h11;
assign _c_characterGenerator[2819] = 8'h44;
assign _c_characterGenerator[2820] = 8'h11;
assign _c_characterGenerator[2821] = 8'h44;
assign _c_characterGenerator[2822] = 8'h11;
assign _c_characterGenerator[2823] = 8'h44;
assign _c_characterGenerator[2824] = 8'h11;
assign _c_characterGenerator[2825] = 8'h44;
assign _c_characterGenerator[2826] = 8'h11;
assign _c_characterGenerator[2827] = 8'h44;
assign _c_characterGenerator[2828] = 8'h11;
assign _c_characterGenerator[2829] = 8'h44;
assign _c_characterGenerator[2830] = 8'h11;
assign _c_characterGenerator[2831] = 8'h44;
assign _c_characterGenerator[2832] = 8'h55;
assign _c_characterGenerator[2833] = 8'haa;
assign _c_characterGenerator[2834] = 8'h55;
assign _c_characterGenerator[2835] = 8'haa;
assign _c_characterGenerator[2836] = 8'h55;
assign _c_characterGenerator[2837] = 8'haa;
assign _c_characterGenerator[2838] = 8'h55;
assign _c_characterGenerator[2839] = 8'haa;
assign _c_characterGenerator[2840] = 8'h55;
assign _c_characterGenerator[2841] = 8'haa;
assign _c_characterGenerator[2842] = 8'h55;
assign _c_characterGenerator[2843] = 8'haa;
assign _c_characterGenerator[2844] = 8'h55;
assign _c_characterGenerator[2845] = 8'haa;
assign _c_characterGenerator[2846] = 8'h55;
assign _c_characterGenerator[2847] = 8'haa;
assign _c_characterGenerator[2848] = 8'hdd;
assign _c_characterGenerator[2849] = 8'h77;
assign _c_characterGenerator[2850] = 8'hdd;
assign _c_characterGenerator[2851] = 8'h77;
assign _c_characterGenerator[2852] = 8'hdd;
assign _c_characterGenerator[2853] = 8'h77;
assign _c_characterGenerator[2854] = 8'hdd;
assign _c_characterGenerator[2855] = 8'h77;
assign _c_characterGenerator[2856] = 8'hdd;
assign _c_characterGenerator[2857] = 8'h77;
assign _c_characterGenerator[2858] = 8'hdd;
assign _c_characterGenerator[2859] = 8'h77;
assign _c_characterGenerator[2860] = 8'hdd;
assign _c_characterGenerator[2861] = 8'h77;
assign _c_characterGenerator[2862] = 8'hdd;
assign _c_characterGenerator[2863] = 8'h77;
assign _c_characterGenerator[2864] = 8'h18;
assign _c_characterGenerator[2865] = 8'h18;
assign _c_characterGenerator[2866] = 8'h18;
assign _c_characterGenerator[2867] = 8'h18;
assign _c_characterGenerator[2868] = 8'h18;
assign _c_characterGenerator[2869] = 8'h18;
assign _c_characterGenerator[2870] = 8'h18;
assign _c_characterGenerator[2871] = 8'h18;
assign _c_characterGenerator[2872] = 8'h18;
assign _c_characterGenerator[2873] = 8'h18;
assign _c_characterGenerator[2874] = 8'h18;
assign _c_characterGenerator[2875] = 8'h18;
assign _c_characterGenerator[2876] = 8'h18;
assign _c_characterGenerator[2877] = 8'h18;
assign _c_characterGenerator[2878] = 8'h18;
assign _c_characterGenerator[2879] = 8'h18;
assign _c_characterGenerator[2880] = 8'h18;
assign _c_characterGenerator[2881] = 8'h18;
assign _c_characterGenerator[2882] = 8'h18;
assign _c_characterGenerator[2883] = 8'h18;
assign _c_characterGenerator[2884] = 8'h18;
assign _c_characterGenerator[2885] = 8'h18;
assign _c_characterGenerator[2886] = 8'h18;
assign _c_characterGenerator[2887] = 8'hf8;
assign _c_characterGenerator[2888] = 8'h18;
assign _c_characterGenerator[2889] = 8'h18;
assign _c_characterGenerator[2890] = 8'h18;
assign _c_characterGenerator[2891] = 8'h18;
assign _c_characterGenerator[2892] = 8'h18;
assign _c_characterGenerator[2893] = 8'h18;
assign _c_characterGenerator[2894] = 8'h18;
assign _c_characterGenerator[2895] = 8'h18;
assign _c_characterGenerator[2896] = 8'h18;
assign _c_characterGenerator[2897] = 8'h18;
assign _c_characterGenerator[2898] = 8'h18;
assign _c_characterGenerator[2899] = 8'h18;
assign _c_characterGenerator[2900] = 8'h18;
assign _c_characterGenerator[2901] = 8'hf8;
assign _c_characterGenerator[2902] = 8'h18;
assign _c_characterGenerator[2903] = 8'hf8;
assign _c_characterGenerator[2904] = 8'h18;
assign _c_characterGenerator[2905] = 8'h18;
assign _c_characterGenerator[2906] = 8'h18;
assign _c_characterGenerator[2907] = 8'h18;
assign _c_characterGenerator[2908] = 8'h18;
assign _c_characterGenerator[2909] = 8'h18;
assign _c_characterGenerator[2910] = 8'h18;
assign _c_characterGenerator[2911] = 8'h18;
assign _c_characterGenerator[2912] = 8'h36;
assign _c_characterGenerator[2913] = 8'h36;
assign _c_characterGenerator[2914] = 8'h36;
assign _c_characterGenerator[2915] = 8'h36;
assign _c_characterGenerator[2916] = 8'h36;
assign _c_characterGenerator[2917] = 8'h36;
assign _c_characterGenerator[2918] = 8'h36;
assign _c_characterGenerator[2919] = 8'hf6;
assign _c_characterGenerator[2920] = 8'h36;
assign _c_characterGenerator[2921] = 8'h36;
assign _c_characterGenerator[2922] = 8'h36;
assign _c_characterGenerator[2923] = 8'h36;
assign _c_characterGenerator[2924] = 8'h36;
assign _c_characterGenerator[2925] = 8'h36;
assign _c_characterGenerator[2926] = 8'h36;
assign _c_characterGenerator[2927] = 8'h36;
assign _c_characterGenerator[2928] = 8'h00;
assign _c_characterGenerator[2929] = 8'h00;
assign _c_characterGenerator[2930] = 8'h00;
assign _c_characterGenerator[2931] = 8'h00;
assign _c_characterGenerator[2932] = 8'h00;
assign _c_characterGenerator[2933] = 8'h00;
assign _c_characterGenerator[2934] = 8'h00;
assign _c_characterGenerator[2935] = 8'hfe;
assign _c_characterGenerator[2936] = 8'h36;
assign _c_characterGenerator[2937] = 8'h36;
assign _c_characterGenerator[2938] = 8'h36;
assign _c_characterGenerator[2939] = 8'h36;
assign _c_characterGenerator[2940] = 8'h36;
assign _c_characterGenerator[2941] = 8'h36;
assign _c_characterGenerator[2942] = 8'h36;
assign _c_characterGenerator[2943] = 8'h36;
assign _c_characterGenerator[2944] = 8'h00;
assign _c_characterGenerator[2945] = 8'h00;
assign _c_characterGenerator[2946] = 8'h00;
assign _c_characterGenerator[2947] = 8'h00;
assign _c_characterGenerator[2948] = 8'h00;
assign _c_characterGenerator[2949] = 8'hf8;
assign _c_characterGenerator[2950] = 8'h18;
assign _c_characterGenerator[2951] = 8'hf8;
assign _c_characterGenerator[2952] = 8'h18;
assign _c_characterGenerator[2953] = 8'h18;
assign _c_characterGenerator[2954] = 8'h18;
assign _c_characterGenerator[2955] = 8'h18;
assign _c_characterGenerator[2956] = 8'h18;
assign _c_characterGenerator[2957] = 8'h18;
assign _c_characterGenerator[2958] = 8'h18;
assign _c_characterGenerator[2959] = 8'h18;
assign _c_characterGenerator[2960] = 8'h36;
assign _c_characterGenerator[2961] = 8'h36;
assign _c_characterGenerator[2962] = 8'h36;
assign _c_characterGenerator[2963] = 8'h36;
assign _c_characterGenerator[2964] = 8'h36;
assign _c_characterGenerator[2965] = 8'hf6;
assign _c_characterGenerator[2966] = 8'h06;
assign _c_characterGenerator[2967] = 8'hf6;
assign _c_characterGenerator[2968] = 8'h36;
assign _c_characterGenerator[2969] = 8'h36;
assign _c_characterGenerator[2970] = 8'h36;
assign _c_characterGenerator[2971] = 8'h36;
assign _c_characterGenerator[2972] = 8'h36;
assign _c_characterGenerator[2973] = 8'h36;
assign _c_characterGenerator[2974] = 8'h36;
assign _c_characterGenerator[2975] = 8'h36;
assign _c_characterGenerator[2976] = 8'h36;
assign _c_characterGenerator[2977] = 8'h36;
assign _c_characterGenerator[2978] = 8'h36;
assign _c_characterGenerator[2979] = 8'h36;
assign _c_characterGenerator[2980] = 8'h36;
assign _c_characterGenerator[2981] = 8'h36;
assign _c_characterGenerator[2982] = 8'h36;
assign _c_characterGenerator[2983] = 8'h36;
assign _c_characterGenerator[2984] = 8'h36;
assign _c_characterGenerator[2985] = 8'h36;
assign _c_characterGenerator[2986] = 8'h36;
assign _c_characterGenerator[2987] = 8'h36;
assign _c_characterGenerator[2988] = 8'h36;
assign _c_characterGenerator[2989] = 8'h36;
assign _c_characterGenerator[2990] = 8'h36;
assign _c_characterGenerator[2991] = 8'h36;
assign _c_characterGenerator[2992] = 8'h00;
assign _c_characterGenerator[2993] = 8'h00;
assign _c_characterGenerator[2994] = 8'h00;
assign _c_characterGenerator[2995] = 8'h00;
assign _c_characterGenerator[2996] = 8'h00;
assign _c_characterGenerator[2997] = 8'hfe;
assign _c_characterGenerator[2998] = 8'h06;
assign _c_characterGenerator[2999] = 8'hf6;
assign _c_characterGenerator[3000] = 8'h36;
assign _c_characterGenerator[3001] = 8'h36;
assign _c_characterGenerator[3002] = 8'h36;
assign _c_characterGenerator[3003] = 8'h36;
assign _c_characterGenerator[3004] = 8'h36;
assign _c_characterGenerator[3005] = 8'h36;
assign _c_characterGenerator[3006] = 8'h36;
assign _c_characterGenerator[3007] = 8'h36;
assign _c_characterGenerator[3008] = 8'h36;
assign _c_characterGenerator[3009] = 8'h36;
assign _c_characterGenerator[3010] = 8'h36;
assign _c_characterGenerator[3011] = 8'h36;
assign _c_characterGenerator[3012] = 8'h36;
assign _c_characterGenerator[3013] = 8'hf6;
assign _c_characterGenerator[3014] = 8'h06;
assign _c_characterGenerator[3015] = 8'hfe;
assign _c_characterGenerator[3016] = 8'h00;
assign _c_characterGenerator[3017] = 8'h00;
assign _c_characterGenerator[3018] = 8'h00;
assign _c_characterGenerator[3019] = 8'h00;
assign _c_characterGenerator[3020] = 8'h00;
assign _c_characterGenerator[3021] = 8'h00;
assign _c_characterGenerator[3022] = 8'h00;
assign _c_characterGenerator[3023] = 8'h00;
assign _c_characterGenerator[3024] = 8'h36;
assign _c_characterGenerator[3025] = 8'h36;
assign _c_characterGenerator[3026] = 8'h36;
assign _c_characterGenerator[3027] = 8'h36;
assign _c_characterGenerator[3028] = 8'h36;
assign _c_characterGenerator[3029] = 8'h36;
assign _c_characterGenerator[3030] = 8'h36;
assign _c_characterGenerator[3031] = 8'hfe;
assign _c_characterGenerator[3032] = 8'h00;
assign _c_characterGenerator[3033] = 8'h00;
assign _c_characterGenerator[3034] = 8'h00;
assign _c_characterGenerator[3035] = 8'h00;
assign _c_characterGenerator[3036] = 8'h00;
assign _c_characterGenerator[3037] = 8'h00;
assign _c_characterGenerator[3038] = 8'h00;
assign _c_characterGenerator[3039] = 8'h00;
assign _c_characterGenerator[3040] = 8'h18;
assign _c_characterGenerator[3041] = 8'h18;
assign _c_characterGenerator[3042] = 8'h18;
assign _c_characterGenerator[3043] = 8'h18;
assign _c_characterGenerator[3044] = 8'h18;
assign _c_characterGenerator[3045] = 8'hf8;
assign _c_characterGenerator[3046] = 8'h18;
assign _c_characterGenerator[3047] = 8'hf8;
assign _c_characterGenerator[3048] = 8'h00;
assign _c_characterGenerator[3049] = 8'h00;
assign _c_characterGenerator[3050] = 8'h00;
assign _c_characterGenerator[3051] = 8'h00;
assign _c_characterGenerator[3052] = 8'h00;
assign _c_characterGenerator[3053] = 8'h00;
assign _c_characterGenerator[3054] = 8'h00;
assign _c_characterGenerator[3055] = 8'h00;
assign _c_characterGenerator[3056] = 8'h00;
assign _c_characterGenerator[3057] = 8'h00;
assign _c_characterGenerator[3058] = 8'h00;
assign _c_characterGenerator[3059] = 8'h00;
assign _c_characterGenerator[3060] = 8'h00;
assign _c_characterGenerator[3061] = 8'h00;
assign _c_characterGenerator[3062] = 8'h00;
assign _c_characterGenerator[3063] = 8'hf8;
assign _c_characterGenerator[3064] = 8'h18;
assign _c_characterGenerator[3065] = 8'h18;
assign _c_characterGenerator[3066] = 8'h18;
assign _c_characterGenerator[3067] = 8'h18;
assign _c_characterGenerator[3068] = 8'h18;
assign _c_characterGenerator[3069] = 8'h18;
assign _c_characterGenerator[3070] = 8'h18;
assign _c_characterGenerator[3071] = 8'h18;
assign _c_characterGenerator[3072] = 8'h18;
assign _c_characterGenerator[3073] = 8'h18;
assign _c_characterGenerator[3074] = 8'h18;
assign _c_characterGenerator[3075] = 8'h18;
assign _c_characterGenerator[3076] = 8'h18;
assign _c_characterGenerator[3077] = 8'h18;
assign _c_characterGenerator[3078] = 8'h18;
assign _c_characterGenerator[3079] = 8'h1f;
assign _c_characterGenerator[3080] = 8'h00;
assign _c_characterGenerator[3081] = 8'h00;
assign _c_characterGenerator[3082] = 8'h00;
assign _c_characterGenerator[3083] = 8'h00;
assign _c_characterGenerator[3084] = 8'h00;
assign _c_characterGenerator[3085] = 8'h00;
assign _c_characterGenerator[3086] = 8'h00;
assign _c_characterGenerator[3087] = 8'h00;
assign _c_characterGenerator[3088] = 8'h18;
assign _c_characterGenerator[3089] = 8'h18;
assign _c_characterGenerator[3090] = 8'h18;
assign _c_characterGenerator[3091] = 8'h18;
assign _c_characterGenerator[3092] = 8'h18;
assign _c_characterGenerator[3093] = 8'h18;
assign _c_characterGenerator[3094] = 8'h18;
assign _c_characterGenerator[3095] = 8'hff;
assign _c_characterGenerator[3096] = 8'h00;
assign _c_characterGenerator[3097] = 8'h00;
assign _c_characterGenerator[3098] = 8'h00;
assign _c_characterGenerator[3099] = 8'h00;
assign _c_characterGenerator[3100] = 8'h00;
assign _c_characterGenerator[3101] = 8'h00;
assign _c_characterGenerator[3102] = 8'h00;
assign _c_characterGenerator[3103] = 8'h00;
assign _c_characterGenerator[3104] = 8'h00;
assign _c_characterGenerator[3105] = 8'h00;
assign _c_characterGenerator[3106] = 8'h00;
assign _c_characterGenerator[3107] = 8'h00;
assign _c_characterGenerator[3108] = 8'h00;
assign _c_characterGenerator[3109] = 8'h00;
assign _c_characterGenerator[3110] = 8'h00;
assign _c_characterGenerator[3111] = 8'hff;
assign _c_characterGenerator[3112] = 8'h18;
assign _c_characterGenerator[3113] = 8'h18;
assign _c_characterGenerator[3114] = 8'h18;
assign _c_characterGenerator[3115] = 8'h18;
assign _c_characterGenerator[3116] = 8'h18;
assign _c_characterGenerator[3117] = 8'h18;
assign _c_characterGenerator[3118] = 8'h18;
assign _c_characterGenerator[3119] = 8'h18;
assign _c_characterGenerator[3120] = 8'h18;
assign _c_characterGenerator[3121] = 8'h18;
assign _c_characterGenerator[3122] = 8'h18;
assign _c_characterGenerator[3123] = 8'h18;
assign _c_characterGenerator[3124] = 8'h18;
assign _c_characterGenerator[3125] = 8'h18;
assign _c_characterGenerator[3126] = 8'h18;
assign _c_characterGenerator[3127] = 8'h1f;
assign _c_characterGenerator[3128] = 8'h18;
assign _c_characterGenerator[3129] = 8'h18;
assign _c_characterGenerator[3130] = 8'h18;
assign _c_characterGenerator[3131] = 8'h18;
assign _c_characterGenerator[3132] = 8'h18;
assign _c_characterGenerator[3133] = 8'h18;
assign _c_characterGenerator[3134] = 8'h18;
assign _c_characterGenerator[3135] = 8'h18;
assign _c_characterGenerator[3136] = 8'h00;
assign _c_characterGenerator[3137] = 8'h00;
assign _c_characterGenerator[3138] = 8'h00;
assign _c_characterGenerator[3139] = 8'h00;
assign _c_characterGenerator[3140] = 8'h00;
assign _c_characterGenerator[3141] = 8'h00;
assign _c_characterGenerator[3142] = 8'h00;
assign _c_characterGenerator[3143] = 8'hff;
assign _c_characterGenerator[3144] = 8'h00;
assign _c_characterGenerator[3145] = 8'h00;
assign _c_characterGenerator[3146] = 8'h00;
assign _c_characterGenerator[3147] = 8'h00;
assign _c_characterGenerator[3148] = 8'h00;
assign _c_characterGenerator[3149] = 8'h00;
assign _c_characterGenerator[3150] = 8'h00;
assign _c_characterGenerator[3151] = 8'h00;
assign _c_characterGenerator[3152] = 8'h18;
assign _c_characterGenerator[3153] = 8'h18;
assign _c_characterGenerator[3154] = 8'h18;
assign _c_characterGenerator[3155] = 8'h18;
assign _c_characterGenerator[3156] = 8'h18;
assign _c_characterGenerator[3157] = 8'h18;
assign _c_characterGenerator[3158] = 8'h18;
assign _c_characterGenerator[3159] = 8'hff;
assign _c_characterGenerator[3160] = 8'h18;
assign _c_characterGenerator[3161] = 8'h18;
assign _c_characterGenerator[3162] = 8'h18;
assign _c_characterGenerator[3163] = 8'h18;
assign _c_characterGenerator[3164] = 8'h18;
assign _c_characterGenerator[3165] = 8'h18;
assign _c_characterGenerator[3166] = 8'h18;
assign _c_characterGenerator[3167] = 8'h18;
assign _c_characterGenerator[3168] = 8'h18;
assign _c_characterGenerator[3169] = 8'h18;
assign _c_characterGenerator[3170] = 8'h18;
assign _c_characterGenerator[3171] = 8'h18;
assign _c_characterGenerator[3172] = 8'h18;
assign _c_characterGenerator[3173] = 8'h1f;
assign _c_characterGenerator[3174] = 8'h18;
assign _c_characterGenerator[3175] = 8'h1f;
assign _c_characterGenerator[3176] = 8'h18;
assign _c_characterGenerator[3177] = 8'h18;
assign _c_characterGenerator[3178] = 8'h18;
assign _c_characterGenerator[3179] = 8'h18;
assign _c_characterGenerator[3180] = 8'h18;
assign _c_characterGenerator[3181] = 8'h18;
assign _c_characterGenerator[3182] = 8'h18;
assign _c_characterGenerator[3183] = 8'h18;
assign _c_characterGenerator[3184] = 8'h36;
assign _c_characterGenerator[3185] = 8'h36;
assign _c_characterGenerator[3186] = 8'h36;
assign _c_characterGenerator[3187] = 8'h36;
assign _c_characterGenerator[3188] = 8'h36;
assign _c_characterGenerator[3189] = 8'h36;
assign _c_characterGenerator[3190] = 8'h36;
assign _c_characterGenerator[3191] = 8'h37;
assign _c_characterGenerator[3192] = 8'h36;
assign _c_characterGenerator[3193] = 8'h36;
assign _c_characterGenerator[3194] = 8'h36;
assign _c_characterGenerator[3195] = 8'h36;
assign _c_characterGenerator[3196] = 8'h36;
assign _c_characterGenerator[3197] = 8'h36;
assign _c_characterGenerator[3198] = 8'h36;
assign _c_characterGenerator[3199] = 8'h36;
assign _c_characterGenerator[3200] = 8'h36;
assign _c_characterGenerator[3201] = 8'h36;
assign _c_characterGenerator[3202] = 8'h36;
assign _c_characterGenerator[3203] = 8'h36;
assign _c_characterGenerator[3204] = 8'h36;
assign _c_characterGenerator[3205] = 8'h37;
assign _c_characterGenerator[3206] = 8'h30;
assign _c_characterGenerator[3207] = 8'h3f;
assign _c_characterGenerator[3208] = 8'h00;
assign _c_characterGenerator[3209] = 8'h00;
assign _c_characterGenerator[3210] = 8'h00;
assign _c_characterGenerator[3211] = 8'h00;
assign _c_characterGenerator[3212] = 8'h00;
assign _c_characterGenerator[3213] = 8'h00;
assign _c_characterGenerator[3214] = 8'h00;
assign _c_characterGenerator[3215] = 8'h00;
assign _c_characterGenerator[3216] = 8'h00;
assign _c_characterGenerator[3217] = 8'h00;
assign _c_characterGenerator[3218] = 8'h00;
assign _c_characterGenerator[3219] = 8'h00;
assign _c_characterGenerator[3220] = 8'h00;
assign _c_characterGenerator[3221] = 8'h3f;
assign _c_characterGenerator[3222] = 8'h30;
assign _c_characterGenerator[3223] = 8'h37;
assign _c_characterGenerator[3224] = 8'h36;
assign _c_characterGenerator[3225] = 8'h36;
assign _c_characterGenerator[3226] = 8'h36;
assign _c_characterGenerator[3227] = 8'h36;
assign _c_characterGenerator[3228] = 8'h36;
assign _c_characterGenerator[3229] = 8'h36;
assign _c_characterGenerator[3230] = 8'h36;
assign _c_characterGenerator[3231] = 8'h36;
assign _c_characterGenerator[3232] = 8'h36;
assign _c_characterGenerator[3233] = 8'h36;
assign _c_characterGenerator[3234] = 8'h36;
assign _c_characterGenerator[3235] = 8'h36;
assign _c_characterGenerator[3236] = 8'h36;
assign _c_characterGenerator[3237] = 8'hf7;
assign _c_characterGenerator[3238] = 8'h00;
assign _c_characterGenerator[3239] = 8'hff;
assign _c_characterGenerator[3240] = 8'h00;
assign _c_characterGenerator[3241] = 8'h00;
assign _c_characterGenerator[3242] = 8'h00;
assign _c_characterGenerator[3243] = 8'h00;
assign _c_characterGenerator[3244] = 8'h00;
assign _c_characterGenerator[3245] = 8'h00;
assign _c_characterGenerator[3246] = 8'h00;
assign _c_characterGenerator[3247] = 8'h00;
assign _c_characterGenerator[3248] = 8'h00;
assign _c_characterGenerator[3249] = 8'h00;
assign _c_characterGenerator[3250] = 8'h00;
assign _c_characterGenerator[3251] = 8'h00;
assign _c_characterGenerator[3252] = 8'h00;
assign _c_characterGenerator[3253] = 8'hff;
assign _c_characterGenerator[3254] = 8'h00;
assign _c_characterGenerator[3255] = 8'hf7;
assign _c_characterGenerator[3256] = 8'h36;
assign _c_characterGenerator[3257] = 8'h36;
assign _c_characterGenerator[3258] = 8'h36;
assign _c_characterGenerator[3259] = 8'h36;
assign _c_characterGenerator[3260] = 8'h36;
assign _c_characterGenerator[3261] = 8'h36;
assign _c_characterGenerator[3262] = 8'h36;
assign _c_characterGenerator[3263] = 8'h36;
assign _c_characterGenerator[3264] = 8'h36;
assign _c_characterGenerator[3265] = 8'h36;
assign _c_characterGenerator[3266] = 8'h36;
assign _c_characterGenerator[3267] = 8'h36;
assign _c_characterGenerator[3268] = 8'h36;
assign _c_characterGenerator[3269] = 8'h37;
assign _c_characterGenerator[3270] = 8'h30;
assign _c_characterGenerator[3271] = 8'h37;
assign _c_characterGenerator[3272] = 8'h36;
assign _c_characterGenerator[3273] = 8'h36;
assign _c_characterGenerator[3274] = 8'h36;
assign _c_characterGenerator[3275] = 8'h36;
assign _c_characterGenerator[3276] = 8'h36;
assign _c_characterGenerator[3277] = 8'h36;
assign _c_characterGenerator[3278] = 8'h36;
assign _c_characterGenerator[3279] = 8'h36;
assign _c_characterGenerator[3280] = 8'h00;
assign _c_characterGenerator[3281] = 8'h00;
assign _c_characterGenerator[3282] = 8'h00;
assign _c_characterGenerator[3283] = 8'h00;
assign _c_characterGenerator[3284] = 8'h00;
assign _c_characterGenerator[3285] = 8'hff;
assign _c_characterGenerator[3286] = 8'h00;
assign _c_characterGenerator[3287] = 8'hff;
assign _c_characterGenerator[3288] = 8'h00;
assign _c_characterGenerator[3289] = 8'h00;
assign _c_characterGenerator[3290] = 8'h00;
assign _c_characterGenerator[3291] = 8'h00;
assign _c_characterGenerator[3292] = 8'h00;
assign _c_characterGenerator[3293] = 8'h00;
assign _c_characterGenerator[3294] = 8'h00;
assign _c_characterGenerator[3295] = 8'h00;
assign _c_characterGenerator[3296] = 8'h36;
assign _c_characterGenerator[3297] = 8'h36;
assign _c_characterGenerator[3298] = 8'h36;
assign _c_characterGenerator[3299] = 8'h36;
assign _c_characterGenerator[3300] = 8'h36;
assign _c_characterGenerator[3301] = 8'hf7;
assign _c_characterGenerator[3302] = 8'h00;
assign _c_characterGenerator[3303] = 8'hf7;
assign _c_characterGenerator[3304] = 8'h36;
assign _c_characterGenerator[3305] = 8'h36;
assign _c_characterGenerator[3306] = 8'h36;
assign _c_characterGenerator[3307] = 8'h36;
assign _c_characterGenerator[3308] = 8'h36;
assign _c_characterGenerator[3309] = 8'h36;
assign _c_characterGenerator[3310] = 8'h36;
assign _c_characterGenerator[3311] = 8'h36;
assign _c_characterGenerator[3312] = 8'h18;
assign _c_characterGenerator[3313] = 8'h18;
assign _c_characterGenerator[3314] = 8'h18;
assign _c_characterGenerator[3315] = 8'h18;
assign _c_characterGenerator[3316] = 8'h18;
assign _c_characterGenerator[3317] = 8'hff;
assign _c_characterGenerator[3318] = 8'h00;
assign _c_characterGenerator[3319] = 8'hff;
assign _c_characterGenerator[3320] = 8'h00;
assign _c_characterGenerator[3321] = 8'h00;
assign _c_characterGenerator[3322] = 8'h00;
assign _c_characterGenerator[3323] = 8'h00;
assign _c_characterGenerator[3324] = 8'h00;
assign _c_characterGenerator[3325] = 8'h00;
assign _c_characterGenerator[3326] = 8'h00;
assign _c_characterGenerator[3327] = 8'h00;
assign _c_characterGenerator[3328] = 8'h36;
assign _c_characterGenerator[3329] = 8'h36;
assign _c_characterGenerator[3330] = 8'h36;
assign _c_characterGenerator[3331] = 8'h36;
assign _c_characterGenerator[3332] = 8'h36;
assign _c_characterGenerator[3333] = 8'h36;
assign _c_characterGenerator[3334] = 8'h36;
assign _c_characterGenerator[3335] = 8'hff;
assign _c_characterGenerator[3336] = 8'h00;
assign _c_characterGenerator[3337] = 8'h00;
assign _c_characterGenerator[3338] = 8'h00;
assign _c_characterGenerator[3339] = 8'h00;
assign _c_characterGenerator[3340] = 8'h00;
assign _c_characterGenerator[3341] = 8'h00;
assign _c_characterGenerator[3342] = 8'h00;
assign _c_characterGenerator[3343] = 8'h00;
assign _c_characterGenerator[3344] = 8'h00;
assign _c_characterGenerator[3345] = 8'h00;
assign _c_characterGenerator[3346] = 8'h00;
assign _c_characterGenerator[3347] = 8'h00;
assign _c_characterGenerator[3348] = 8'h00;
assign _c_characterGenerator[3349] = 8'hff;
assign _c_characterGenerator[3350] = 8'h00;
assign _c_characterGenerator[3351] = 8'hff;
assign _c_characterGenerator[3352] = 8'h18;
assign _c_characterGenerator[3353] = 8'h18;
assign _c_characterGenerator[3354] = 8'h18;
assign _c_characterGenerator[3355] = 8'h18;
assign _c_characterGenerator[3356] = 8'h18;
assign _c_characterGenerator[3357] = 8'h18;
assign _c_characterGenerator[3358] = 8'h18;
assign _c_characterGenerator[3359] = 8'h18;
assign _c_characterGenerator[3360] = 8'h00;
assign _c_characterGenerator[3361] = 8'h00;
assign _c_characterGenerator[3362] = 8'h00;
assign _c_characterGenerator[3363] = 8'h00;
assign _c_characterGenerator[3364] = 8'h00;
assign _c_characterGenerator[3365] = 8'h00;
assign _c_characterGenerator[3366] = 8'h00;
assign _c_characterGenerator[3367] = 8'hff;
assign _c_characterGenerator[3368] = 8'h36;
assign _c_characterGenerator[3369] = 8'h36;
assign _c_characterGenerator[3370] = 8'h36;
assign _c_characterGenerator[3371] = 8'h36;
assign _c_characterGenerator[3372] = 8'h36;
assign _c_characterGenerator[3373] = 8'h36;
assign _c_characterGenerator[3374] = 8'h36;
assign _c_characterGenerator[3375] = 8'h36;
assign _c_characterGenerator[3376] = 8'h36;
assign _c_characterGenerator[3377] = 8'h36;
assign _c_characterGenerator[3378] = 8'h36;
assign _c_characterGenerator[3379] = 8'h36;
assign _c_characterGenerator[3380] = 8'h36;
assign _c_characterGenerator[3381] = 8'h36;
assign _c_characterGenerator[3382] = 8'h36;
assign _c_characterGenerator[3383] = 8'h3f;
assign _c_characterGenerator[3384] = 8'h00;
assign _c_characterGenerator[3385] = 8'h00;
assign _c_characterGenerator[3386] = 8'h00;
assign _c_characterGenerator[3387] = 8'h00;
assign _c_characterGenerator[3388] = 8'h00;
assign _c_characterGenerator[3389] = 8'h00;
assign _c_characterGenerator[3390] = 8'h00;
assign _c_characterGenerator[3391] = 8'h00;
assign _c_characterGenerator[3392] = 8'h18;
assign _c_characterGenerator[3393] = 8'h18;
assign _c_characterGenerator[3394] = 8'h18;
assign _c_characterGenerator[3395] = 8'h18;
assign _c_characterGenerator[3396] = 8'h18;
assign _c_characterGenerator[3397] = 8'h1f;
assign _c_characterGenerator[3398] = 8'h18;
assign _c_characterGenerator[3399] = 8'h1f;
assign _c_characterGenerator[3400] = 8'h00;
assign _c_characterGenerator[3401] = 8'h00;
assign _c_characterGenerator[3402] = 8'h00;
assign _c_characterGenerator[3403] = 8'h00;
assign _c_characterGenerator[3404] = 8'h00;
assign _c_characterGenerator[3405] = 8'h00;
assign _c_characterGenerator[3406] = 8'h00;
assign _c_characterGenerator[3407] = 8'h00;
assign _c_characterGenerator[3408] = 8'h00;
assign _c_characterGenerator[3409] = 8'h00;
assign _c_characterGenerator[3410] = 8'h00;
assign _c_characterGenerator[3411] = 8'h00;
assign _c_characterGenerator[3412] = 8'h00;
assign _c_characterGenerator[3413] = 8'h1f;
assign _c_characterGenerator[3414] = 8'h18;
assign _c_characterGenerator[3415] = 8'h1f;
assign _c_characterGenerator[3416] = 8'h18;
assign _c_characterGenerator[3417] = 8'h18;
assign _c_characterGenerator[3418] = 8'h18;
assign _c_characterGenerator[3419] = 8'h18;
assign _c_characterGenerator[3420] = 8'h18;
assign _c_characterGenerator[3421] = 8'h18;
assign _c_characterGenerator[3422] = 8'h18;
assign _c_characterGenerator[3423] = 8'h18;
assign _c_characterGenerator[3424] = 8'h00;
assign _c_characterGenerator[3425] = 8'h00;
assign _c_characterGenerator[3426] = 8'h00;
assign _c_characterGenerator[3427] = 8'h00;
assign _c_characterGenerator[3428] = 8'h00;
assign _c_characterGenerator[3429] = 8'h00;
assign _c_characterGenerator[3430] = 8'h00;
assign _c_characterGenerator[3431] = 8'h3f;
assign _c_characterGenerator[3432] = 8'h36;
assign _c_characterGenerator[3433] = 8'h36;
assign _c_characterGenerator[3434] = 8'h36;
assign _c_characterGenerator[3435] = 8'h36;
assign _c_characterGenerator[3436] = 8'h36;
assign _c_characterGenerator[3437] = 8'h36;
assign _c_characterGenerator[3438] = 8'h36;
assign _c_characterGenerator[3439] = 8'h36;
assign _c_characterGenerator[3440] = 8'h36;
assign _c_characterGenerator[3441] = 8'h36;
assign _c_characterGenerator[3442] = 8'h36;
assign _c_characterGenerator[3443] = 8'h36;
assign _c_characterGenerator[3444] = 8'h36;
assign _c_characterGenerator[3445] = 8'h36;
assign _c_characterGenerator[3446] = 8'h36;
assign _c_characterGenerator[3447] = 8'hff;
assign _c_characterGenerator[3448] = 8'h36;
assign _c_characterGenerator[3449] = 8'h36;
assign _c_characterGenerator[3450] = 8'h36;
assign _c_characterGenerator[3451] = 8'h36;
assign _c_characterGenerator[3452] = 8'h36;
assign _c_characterGenerator[3453] = 8'h36;
assign _c_characterGenerator[3454] = 8'h36;
assign _c_characterGenerator[3455] = 8'h36;
assign _c_characterGenerator[3456] = 8'h18;
assign _c_characterGenerator[3457] = 8'h18;
assign _c_characterGenerator[3458] = 8'h18;
assign _c_characterGenerator[3459] = 8'h18;
assign _c_characterGenerator[3460] = 8'h18;
assign _c_characterGenerator[3461] = 8'hff;
assign _c_characterGenerator[3462] = 8'h18;
assign _c_characterGenerator[3463] = 8'hff;
assign _c_characterGenerator[3464] = 8'h18;
assign _c_characterGenerator[3465] = 8'h18;
assign _c_characterGenerator[3466] = 8'h18;
assign _c_characterGenerator[3467] = 8'h18;
assign _c_characterGenerator[3468] = 8'h18;
assign _c_characterGenerator[3469] = 8'h18;
assign _c_characterGenerator[3470] = 8'h18;
assign _c_characterGenerator[3471] = 8'h18;
assign _c_characterGenerator[3472] = 8'h18;
assign _c_characterGenerator[3473] = 8'h18;
assign _c_characterGenerator[3474] = 8'h18;
assign _c_characterGenerator[3475] = 8'h18;
assign _c_characterGenerator[3476] = 8'h18;
assign _c_characterGenerator[3477] = 8'h18;
assign _c_characterGenerator[3478] = 8'h18;
assign _c_characterGenerator[3479] = 8'hf8;
assign _c_characterGenerator[3480] = 8'h00;
assign _c_characterGenerator[3481] = 8'h00;
assign _c_characterGenerator[3482] = 8'h00;
assign _c_characterGenerator[3483] = 8'h00;
assign _c_characterGenerator[3484] = 8'h00;
assign _c_characterGenerator[3485] = 8'h00;
assign _c_characterGenerator[3486] = 8'h00;
assign _c_characterGenerator[3487] = 8'h00;
assign _c_characterGenerator[3488] = 8'h00;
assign _c_characterGenerator[3489] = 8'h00;
assign _c_characterGenerator[3490] = 8'h00;
assign _c_characterGenerator[3491] = 8'h00;
assign _c_characterGenerator[3492] = 8'h00;
assign _c_characterGenerator[3493] = 8'h00;
assign _c_characterGenerator[3494] = 8'h00;
assign _c_characterGenerator[3495] = 8'h1f;
assign _c_characterGenerator[3496] = 8'h18;
assign _c_characterGenerator[3497] = 8'h18;
assign _c_characterGenerator[3498] = 8'h18;
assign _c_characterGenerator[3499] = 8'h18;
assign _c_characterGenerator[3500] = 8'h18;
assign _c_characterGenerator[3501] = 8'h18;
assign _c_characterGenerator[3502] = 8'h18;
assign _c_characterGenerator[3503] = 8'h18;
assign _c_characterGenerator[3504] = 8'hff;
assign _c_characterGenerator[3505] = 8'hff;
assign _c_characterGenerator[3506] = 8'hff;
assign _c_characterGenerator[3507] = 8'hff;
assign _c_characterGenerator[3508] = 8'hff;
assign _c_characterGenerator[3509] = 8'hff;
assign _c_characterGenerator[3510] = 8'hff;
assign _c_characterGenerator[3511] = 8'hff;
assign _c_characterGenerator[3512] = 8'hff;
assign _c_characterGenerator[3513] = 8'hff;
assign _c_characterGenerator[3514] = 8'hff;
assign _c_characterGenerator[3515] = 8'hff;
assign _c_characterGenerator[3516] = 8'hff;
assign _c_characterGenerator[3517] = 8'hff;
assign _c_characterGenerator[3518] = 8'hff;
assign _c_characterGenerator[3519] = 8'hff;
assign _c_characterGenerator[3520] = 8'h00;
assign _c_characterGenerator[3521] = 8'h00;
assign _c_characterGenerator[3522] = 8'h00;
assign _c_characterGenerator[3523] = 8'h00;
assign _c_characterGenerator[3524] = 8'h00;
assign _c_characterGenerator[3525] = 8'h00;
assign _c_characterGenerator[3526] = 8'h00;
assign _c_characterGenerator[3527] = 8'hff;
assign _c_characterGenerator[3528] = 8'hff;
assign _c_characterGenerator[3529] = 8'hff;
assign _c_characterGenerator[3530] = 8'hff;
assign _c_characterGenerator[3531] = 8'hff;
assign _c_characterGenerator[3532] = 8'hff;
assign _c_characterGenerator[3533] = 8'hff;
assign _c_characterGenerator[3534] = 8'hff;
assign _c_characterGenerator[3535] = 8'hff;
assign _c_characterGenerator[3536] = 8'hf0;
assign _c_characterGenerator[3537] = 8'hf0;
assign _c_characterGenerator[3538] = 8'hf0;
assign _c_characterGenerator[3539] = 8'hf0;
assign _c_characterGenerator[3540] = 8'hf0;
assign _c_characterGenerator[3541] = 8'hf0;
assign _c_characterGenerator[3542] = 8'hf0;
assign _c_characterGenerator[3543] = 8'hf0;
assign _c_characterGenerator[3544] = 8'hf0;
assign _c_characterGenerator[3545] = 8'hf0;
assign _c_characterGenerator[3546] = 8'hf0;
assign _c_characterGenerator[3547] = 8'hf0;
assign _c_characterGenerator[3548] = 8'hf0;
assign _c_characterGenerator[3549] = 8'hf0;
assign _c_characterGenerator[3550] = 8'hf0;
assign _c_characterGenerator[3551] = 8'hf0;
assign _c_characterGenerator[3552] = 8'h0f;
assign _c_characterGenerator[3553] = 8'h0f;
assign _c_characterGenerator[3554] = 8'h0f;
assign _c_characterGenerator[3555] = 8'h0f;
assign _c_characterGenerator[3556] = 8'h0f;
assign _c_characterGenerator[3557] = 8'h0f;
assign _c_characterGenerator[3558] = 8'h0f;
assign _c_characterGenerator[3559] = 8'h0f;
assign _c_characterGenerator[3560] = 8'h0f;
assign _c_characterGenerator[3561] = 8'h0f;
assign _c_characterGenerator[3562] = 8'h0f;
assign _c_characterGenerator[3563] = 8'h0f;
assign _c_characterGenerator[3564] = 8'h0f;
assign _c_characterGenerator[3565] = 8'h0f;
assign _c_characterGenerator[3566] = 8'h0f;
assign _c_characterGenerator[3567] = 8'h0f;
assign _c_characterGenerator[3568] = 8'hff;
assign _c_characterGenerator[3569] = 8'hff;
assign _c_characterGenerator[3570] = 8'hff;
assign _c_characterGenerator[3571] = 8'hff;
assign _c_characterGenerator[3572] = 8'hff;
assign _c_characterGenerator[3573] = 8'hff;
assign _c_characterGenerator[3574] = 8'hff;
assign _c_characterGenerator[3575] = 8'h00;
assign _c_characterGenerator[3576] = 8'h00;
assign _c_characterGenerator[3577] = 8'h00;
assign _c_characterGenerator[3578] = 8'h00;
assign _c_characterGenerator[3579] = 8'h00;
assign _c_characterGenerator[3580] = 8'h00;
assign _c_characterGenerator[3581] = 8'h00;
assign _c_characterGenerator[3582] = 8'h00;
assign _c_characterGenerator[3583] = 8'h00;
assign _c_characterGenerator[3584] = 8'h00;
assign _c_characterGenerator[3585] = 8'h00;
assign _c_characterGenerator[3586] = 8'h00;
assign _c_characterGenerator[3587] = 8'h00;
assign _c_characterGenerator[3588] = 8'h00;
assign _c_characterGenerator[3589] = 8'h76;
assign _c_characterGenerator[3590] = 8'hdc;
assign _c_characterGenerator[3591] = 8'hd8;
assign _c_characterGenerator[3592] = 8'hd8;
assign _c_characterGenerator[3593] = 8'hd8;
assign _c_characterGenerator[3594] = 8'hdc;
assign _c_characterGenerator[3595] = 8'h76;
assign _c_characterGenerator[3596] = 8'h00;
assign _c_characterGenerator[3597] = 8'h00;
assign _c_characterGenerator[3598] = 8'h00;
assign _c_characterGenerator[3599] = 8'h00;
assign _c_characterGenerator[3600] = 8'h00;
assign _c_characterGenerator[3601] = 8'h00;
assign _c_characterGenerator[3602] = 8'h78;
assign _c_characterGenerator[3603] = 8'hcc;
assign _c_characterGenerator[3604] = 8'hcc;
assign _c_characterGenerator[3605] = 8'hcc;
assign _c_characterGenerator[3606] = 8'hd8;
assign _c_characterGenerator[3607] = 8'hcc;
assign _c_characterGenerator[3608] = 8'hc6;
assign _c_characterGenerator[3609] = 8'hc6;
assign _c_characterGenerator[3610] = 8'hc6;
assign _c_characterGenerator[3611] = 8'hcc;
assign _c_characterGenerator[3612] = 8'h00;
assign _c_characterGenerator[3613] = 8'h00;
assign _c_characterGenerator[3614] = 8'h00;
assign _c_characterGenerator[3615] = 8'h00;
assign _c_characterGenerator[3616] = 8'h00;
assign _c_characterGenerator[3617] = 8'h00;
assign _c_characterGenerator[3618] = 8'hfe;
assign _c_characterGenerator[3619] = 8'hc6;
assign _c_characterGenerator[3620] = 8'hc6;
assign _c_characterGenerator[3621] = 8'hc0;
assign _c_characterGenerator[3622] = 8'hc0;
assign _c_characterGenerator[3623] = 8'hc0;
assign _c_characterGenerator[3624] = 8'hc0;
assign _c_characterGenerator[3625] = 8'hc0;
assign _c_characterGenerator[3626] = 8'hc0;
assign _c_characterGenerator[3627] = 8'hc0;
assign _c_characterGenerator[3628] = 8'h00;
assign _c_characterGenerator[3629] = 8'h00;
assign _c_characterGenerator[3630] = 8'h00;
assign _c_characterGenerator[3631] = 8'h00;
assign _c_characterGenerator[3632] = 8'h00;
assign _c_characterGenerator[3633] = 8'h00;
assign _c_characterGenerator[3634] = 8'h00;
assign _c_characterGenerator[3635] = 8'h00;
assign _c_characterGenerator[3636] = 8'hfe;
assign _c_characterGenerator[3637] = 8'h6c;
assign _c_characterGenerator[3638] = 8'h6c;
assign _c_characterGenerator[3639] = 8'h6c;
assign _c_characterGenerator[3640] = 8'h6c;
assign _c_characterGenerator[3641] = 8'h6c;
assign _c_characterGenerator[3642] = 8'h6c;
assign _c_characterGenerator[3643] = 8'h6c;
assign _c_characterGenerator[3644] = 8'h00;
assign _c_characterGenerator[3645] = 8'h00;
assign _c_characterGenerator[3646] = 8'h00;
assign _c_characterGenerator[3647] = 8'h00;
assign _c_characterGenerator[3648] = 8'h00;
assign _c_characterGenerator[3649] = 8'h00;
assign _c_characterGenerator[3650] = 8'h00;
assign _c_characterGenerator[3651] = 8'hfe;
assign _c_characterGenerator[3652] = 8'hc6;
assign _c_characterGenerator[3653] = 8'h60;
assign _c_characterGenerator[3654] = 8'h30;
assign _c_characterGenerator[3655] = 8'h18;
assign _c_characterGenerator[3656] = 8'h30;
assign _c_characterGenerator[3657] = 8'h60;
assign _c_characterGenerator[3658] = 8'hc6;
assign _c_characterGenerator[3659] = 8'hfe;
assign _c_characterGenerator[3660] = 8'h00;
assign _c_characterGenerator[3661] = 8'h00;
assign _c_characterGenerator[3662] = 8'h00;
assign _c_characterGenerator[3663] = 8'h00;
assign _c_characterGenerator[3664] = 8'h00;
assign _c_characterGenerator[3665] = 8'h00;
assign _c_characterGenerator[3666] = 8'h00;
assign _c_characterGenerator[3667] = 8'h00;
assign _c_characterGenerator[3668] = 8'h00;
assign _c_characterGenerator[3669] = 8'h7e;
assign _c_characterGenerator[3670] = 8'hd8;
assign _c_characterGenerator[3671] = 8'hd8;
assign _c_characterGenerator[3672] = 8'hd8;
assign _c_characterGenerator[3673] = 8'hd8;
assign _c_characterGenerator[3674] = 8'hd8;
assign _c_characterGenerator[3675] = 8'h70;
assign _c_characterGenerator[3676] = 8'h00;
assign _c_characterGenerator[3677] = 8'h00;
assign _c_characterGenerator[3678] = 8'h00;
assign _c_characterGenerator[3679] = 8'h00;
assign _c_characterGenerator[3680] = 8'h00;
assign _c_characterGenerator[3681] = 8'h00;
assign _c_characterGenerator[3682] = 8'h00;
assign _c_characterGenerator[3683] = 8'h00;
assign _c_characterGenerator[3684] = 8'h66;
assign _c_characterGenerator[3685] = 8'h66;
assign _c_characterGenerator[3686] = 8'h66;
assign _c_characterGenerator[3687] = 8'h66;
assign _c_characterGenerator[3688] = 8'h66;
assign _c_characterGenerator[3689] = 8'h7c;
assign _c_characterGenerator[3690] = 8'h60;
assign _c_characterGenerator[3691] = 8'h60;
assign _c_characterGenerator[3692] = 8'hc0;
assign _c_characterGenerator[3693] = 8'h00;
assign _c_characterGenerator[3694] = 8'h00;
assign _c_characterGenerator[3695] = 8'h00;
assign _c_characterGenerator[3696] = 8'h00;
assign _c_characterGenerator[3697] = 8'h00;
assign _c_characterGenerator[3698] = 8'h00;
assign _c_characterGenerator[3699] = 8'h00;
assign _c_characterGenerator[3700] = 8'h76;
assign _c_characterGenerator[3701] = 8'hdc;
assign _c_characterGenerator[3702] = 8'h18;
assign _c_characterGenerator[3703] = 8'h18;
assign _c_characterGenerator[3704] = 8'h18;
assign _c_characterGenerator[3705] = 8'h18;
assign _c_characterGenerator[3706] = 8'h18;
assign _c_characterGenerator[3707] = 8'h18;
assign _c_characterGenerator[3708] = 8'h00;
assign _c_characterGenerator[3709] = 8'h00;
assign _c_characterGenerator[3710] = 8'h00;
assign _c_characterGenerator[3711] = 8'h00;
assign _c_characterGenerator[3712] = 8'h00;
assign _c_characterGenerator[3713] = 8'h00;
assign _c_characterGenerator[3714] = 8'h00;
assign _c_characterGenerator[3715] = 8'h7e;
assign _c_characterGenerator[3716] = 8'h18;
assign _c_characterGenerator[3717] = 8'h3c;
assign _c_characterGenerator[3718] = 8'h66;
assign _c_characterGenerator[3719] = 8'h66;
assign _c_characterGenerator[3720] = 8'h66;
assign _c_characterGenerator[3721] = 8'h3c;
assign _c_characterGenerator[3722] = 8'h18;
assign _c_characterGenerator[3723] = 8'h7e;
assign _c_characterGenerator[3724] = 8'h00;
assign _c_characterGenerator[3725] = 8'h00;
assign _c_characterGenerator[3726] = 8'h00;
assign _c_characterGenerator[3727] = 8'h00;
assign _c_characterGenerator[3728] = 8'h00;
assign _c_characterGenerator[3729] = 8'h00;
assign _c_characterGenerator[3730] = 8'h00;
assign _c_characterGenerator[3731] = 8'h38;
assign _c_characterGenerator[3732] = 8'h6c;
assign _c_characterGenerator[3733] = 8'hc6;
assign _c_characterGenerator[3734] = 8'hc6;
assign _c_characterGenerator[3735] = 8'hfe;
assign _c_characterGenerator[3736] = 8'hc6;
assign _c_characterGenerator[3737] = 8'hc6;
assign _c_characterGenerator[3738] = 8'h6c;
assign _c_characterGenerator[3739] = 8'h38;
assign _c_characterGenerator[3740] = 8'h00;
assign _c_characterGenerator[3741] = 8'h00;
assign _c_characterGenerator[3742] = 8'h00;
assign _c_characterGenerator[3743] = 8'h00;
assign _c_characterGenerator[3744] = 8'h00;
assign _c_characterGenerator[3745] = 8'h00;
assign _c_characterGenerator[3746] = 8'h38;
assign _c_characterGenerator[3747] = 8'h6c;
assign _c_characterGenerator[3748] = 8'hc6;
assign _c_characterGenerator[3749] = 8'hc6;
assign _c_characterGenerator[3750] = 8'hc6;
assign _c_characterGenerator[3751] = 8'h6c;
assign _c_characterGenerator[3752] = 8'h6c;
assign _c_characterGenerator[3753] = 8'h6c;
assign _c_characterGenerator[3754] = 8'h6c;
assign _c_characterGenerator[3755] = 8'hee;
assign _c_characterGenerator[3756] = 8'h00;
assign _c_characterGenerator[3757] = 8'h00;
assign _c_characterGenerator[3758] = 8'h00;
assign _c_characterGenerator[3759] = 8'h00;
assign _c_characterGenerator[3760] = 8'h00;
assign _c_characterGenerator[3761] = 8'h00;
assign _c_characterGenerator[3762] = 8'h1e;
assign _c_characterGenerator[3763] = 8'h30;
assign _c_characterGenerator[3764] = 8'h18;
assign _c_characterGenerator[3765] = 8'h0c;
assign _c_characterGenerator[3766] = 8'h3e;
assign _c_characterGenerator[3767] = 8'h66;
assign _c_characterGenerator[3768] = 8'h66;
assign _c_characterGenerator[3769] = 8'h66;
assign _c_characterGenerator[3770] = 8'h66;
assign _c_characterGenerator[3771] = 8'h3c;
assign _c_characterGenerator[3772] = 8'h00;
assign _c_characterGenerator[3773] = 8'h00;
assign _c_characterGenerator[3774] = 8'h00;
assign _c_characterGenerator[3775] = 8'h00;
assign _c_characterGenerator[3776] = 8'h00;
assign _c_characterGenerator[3777] = 8'h00;
assign _c_characterGenerator[3778] = 8'h00;
assign _c_characterGenerator[3779] = 8'h00;
assign _c_characterGenerator[3780] = 8'h00;
assign _c_characterGenerator[3781] = 8'h7e;
assign _c_characterGenerator[3782] = 8'hdb;
assign _c_characterGenerator[3783] = 8'hdb;
assign _c_characterGenerator[3784] = 8'hdb;
assign _c_characterGenerator[3785] = 8'h7e;
assign _c_characterGenerator[3786] = 8'h00;
assign _c_characterGenerator[3787] = 8'h00;
assign _c_characterGenerator[3788] = 8'h00;
assign _c_characterGenerator[3789] = 8'h00;
assign _c_characterGenerator[3790] = 8'h00;
assign _c_characterGenerator[3791] = 8'h00;
assign _c_characterGenerator[3792] = 8'h00;
assign _c_characterGenerator[3793] = 8'h00;
assign _c_characterGenerator[3794] = 8'h00;
assign _c_characterGenerator[3795] = 8'h03;
assign _c_characterGenerator[3796] = 8'h06;
assign _c_characterGenerator[3797] = 8'h7e;
assign _c_characterGenerator[3798] = 8'hdb;
assign _c_characterGenerator[3799] = 8'hdb;
assign _c_characterGenerator[3800] = 8'hf3;
assign _c_characterGenerator[3801] = 8'h7e;
assign _c_characterGenerator[3802] = 8'h60;
assign _c_characterGenerator[3803] = 8'hc0;
assign _c_characterGenerator[3804] = 8'h00;
assign _c_characterGenerator[3805] = 8'h00;
assign _c_characterGenerator[3806] = 8'h00;
assign _c_characterGenerator[3807] = 8'h00;
assign _c_characterGenerator[3808] = 8'h00;
assign _c_characterGenerator[3809] = 8'h00;
assign _c_characterGenerator[3810] = 8'h1c;
assign _c_characterGenerator[3811] = 8'h30;
assign _c_characterGenerator[3812] = 8'h60;
assign _c_characterGenerator[3813] = 8'h60;
assign _c_characterGenerator[3814] = 8'h7c;
assign _c_characterGenerator[3815] = 8'h60;
assign _c_characterGenerator[3816] = 8'h60;
assign _c_characterGenerator[3817] = 8'h60;
assign _c_characterGenerator[3818] = 8'h30;
assign _c_characterGenerator[3819] = 8'h1c;
assign _c_characterGenerator[3820] = 8'h00;
assign _c_characterGenerator[3821] = 8'h00;
assign _c_characterGenerator[3822] = 8'h00;
assign _c_characterGenerator[3823] = 8'h00;
assign _c_characterGenerator[3824] = 8'h00;
assign _c_characterGenerator[3825] = 8'h00;
assign _c_characterGenerator[3826] = 8'h00;
assign _c_characterGenerator[3827] = 8'h7c;
assign _c_characterGenerator[3828] = 8'hc6;
assign _c_characterGenerator[3829] = 8'hc6;
assign _c_characterGenerator[3830] = 8'hc6;
assign _c_characterGenerator[3831] = 8'hc6;
assign _c_characterGenerator[3832] = 8'hc6;
assign _c_characterGenerator[3833] = 8'hc6;
assign _c_characterGenerator[3834] = 8'hc6;
assign _c_characterGenerator[3835] = 8'hc6;
assign _c_characterGenerator[3836] = 8'h00;
assign _c_characterGenerator[3837] = 8'h00;
assign _c_characterGenerator[3838] = 8'h00;
assign _c_characterGenerator[3839] = 8'h00;
assign _c_characterGenerator[3840] = 8'h00;
assign _c_characterGenerator[3841] = 8'h00;
assign _c_characterGenerator[3842] = 8'h00;
assign _c_characterGenerator[3843] = 8'h00;
assign _c_characterGenerator[3844] = 8'hfe;
assign _c_characterGenerator[3845] = 8'h00;
assign _c_characterGenerator[3846] = 8'h00;
assign _c_characterGenerator[3847] = 8'hfe;
assign _c_characterGenerator[3848] = 8'h00;
assign _c_characterGenerator[3849] = 8'h00;
assign _c_characterGenerator[3850] = 8'hfe;
assign _c_characterGenerator[3851] = 8'h00;
assign _c_characterGenerator[3852] = 8'h00;
assign _c_characterGenerator[3853] = 8'h00;
assign _c_characterGenerator[3854] = 8'h00;
assign _c_characterGenerator[3855] = 8'h00;
assign _c_characterGenerator[3856] = 8'h00;
assign _c_characterGenerator[3857] = 8'h00;
assign _c_characterGenerator[3858] = 8'h00;
assign _c_characterGenerator[3859] = 8'h00;
assign _c_characterGenerator[3860] = 8'h18;
assign _c_characterGenerator[3861] = 8'h18;
assign _c_characterGenerator[3862] = 8'h7e;
assign _c_characterGenerator[3863] = 8'h18;
assign _c_characterGenerator[3864] = 8'h18;
assign _c_characterGenerator[3865] = 8'h00;
assign _c_characterGenerator[3866] = 8'h00;
assign _c_characterGenerator[3867] = 8'hff;
assign _c_characterGenerator[3868] = 8'h00;
assign _c_characterGenerator[3869] = 8'h00;
assign _c_characterGenerator[3870] = 8'h00;
assign _c_characterGenerator[3871] = 8'h00;
assign _c_characterGenerator[3872] = 8'h00;
assign _c_characterGenerator[3873] = 8'h00;
assign _c_characterGenerator[3874] = 8'h00;
assign _c_characterGenerator[3875] = 8'h30;
assign _c_characterGenerator[3876] = 8'h18;
assign _c_characterGenerator[3877] = 8'h0c;
assign _c_characterGenerator[3878] = 8'h06;
assign _c_characterGenerator[3879] = 8'h0c;
assign _c_characterGenerator[3880] = 8'h18;
assign _c_characterGenerator[3881] = 8'h30;
assign _c_characterGenerator[3882] = 8'h00;
assign _c_characterGenerator[3883] = 8'h7e;
assign _c_characterGenerator[3884] = 8'h00;
assign _c_characterGenerator[3885] = 8'h00;
assign _c_characterGenerator[3886] = 8'h00;
assign _c_characterGenerator[3887] = 8'h00;
assign _c_characterGenerator[3888] = 8'h00;
assign _c_characterGenerator[3889] = 8'h00;
assign _c_characterGenerator[3890] = 8'h00;
assign _c_characterGenerator[3891] = 8'h0c;
assign _c_characterGenerator[3892] = 8'h18;
assign _c_characterGenerator[3893] = 8'h30;
assign _c_characterGenerator[3894] = 8'h60;
assign _c_characterGenerator[3895] = 8'h30;
assign _c_characterGenerator[3896] = 8'h18;
assign _c_characterGenerator[3897] = 8'h0c;
assign _c_characterGenerator[3898] = 8'h00;
assign _c_characterGenerator[3899] = 8'h7e;
assign _c_characterGenerator[3900] = 8'h00;
assign _c_characterGenerator[3901] = 8'h00;
assign _c_characterGenerator[3902] = 8'h00;
assign _c_characterGenerator[3903] = 8'h00;
assign _c_characterGenerator[3904] = 8'h00;
assign _c_characterGenerator[3905] = 8'h00;
assign _c_characterGenerator[3906] = 8'h0e;
assign _c_characterGenerator[3907] = 8'h1b;
assign _c_characterGenerator[3908] = 8'h1b;
assign _c_characterGenerator[3909] = 8'h18;
assign _c_characterGenerator[3910] = 8'h18;
assign _c_characterGenerator[3911] = 8'h18;
assign _c_characterGenerator[3912] = 8'h18;
assign _c_characterGenerator[3913] = 8'h18;
assign _c_characterGenerator[3914] = 8'h18;
assign _c_characterGenerator[3915] = 8'h18;
assign _c_characterGenerator[3916] = 8'h18;
assign _c_characterGenerator[3917] = 8'h18;
assign _c_characterGenerator[3918] = 8'h18;
assign _c_characterGenerator[3919] = 8'h18;
assign _c_characterGenerator[3920] = 8'h18;
assign _c_characterGenerator[3921] = 8'h18;
assign _c_characterGenerator[3922] = 8'h18;
assign _c_characterGenerator[3923] = 8'h18;
assign _c_characterGenerator[3924] = 8'h18;
assign _c_characterGenerator[3925] = 8'h18;
assign _c_characterGenerator[3926] = 8'h18;
assign _c_characterGenerator[3927] = 8'h18;
assign _c_characterGenerator[3928] = 8'hd8;
assign _c_characterGenerator[3929] = 8'hd8;
assign _c_characterGenerator[3930] = 8'hd8;
assign _c_characterGenerator[3931] = 8'h70;
assign _c_characterGenerator[3932] = 8'h00;
assign _c_characterGenerator[3933] = 8'h00;
assign _c_characterGenerator[3934] = 8'h00;
assign _c_characterGenerator[3935] = 8'h00;
assign _c_characterGenerator[3936] = 8'h00;
assign _c_characterGenerator[3937] = 8'h00;
assign _c_characterGenerator[3938] = 8'h00;
assign _c_characterGenerator[3939] = 8'h00;
assign _c_characterGenerator[3940] = 8'h18;
assign _c_characterGenerator[3941] = 8'h18;
assign _c_characterGenerator[3942] = 8'h00;
assign _c_characterGenerator[3943] = 8'h7e;
assign _c_characterGenerator[3944] = 8'h00;
assign _c_characterGenerator[3945] = 8'h18;
assign _c_characterGenerator[3946] = 8'h18;
assign _c_characterGenerator[3947] = 8'h00;
assign _c_characterGenerator[3948] = 8'h00;
assign _c_characterGenerator[3949] = 8'h00;
assign _c_characterGenerator[3950] = 8'h00;
assign _c_characterGenerator[3951] = 8'h00;
assign _c_characterGenerator[3952] = 8'h00;
assign _c_characterGenerator[3953] = 8'h00;
assign _c_characterGenerator[3954] = 8'h00;
assign _c_characterGenerator[3955] = 8'h00;
assign _c_characterGenerator[3956] = 8'h00;
assign _c_characterGenerator[3957] = 8'h76;
assign _c_characterGenerator[3958] = 8'hdc;
assign _c_characterGenerator[3959] = 8'h00;
assign _c_characterGenerator[3960] = 8'h76;
assign _c_characterGenerator[3961] = 8'hdc;
assign _c_characterGenerator[3962] = 8'h00;
assign _c_characterGenerator[3963] = 8'h00;
assign _c_characterGenerator[3964] = 8'h00;
assign _c_characterGenerator[3965] = 8'h00;
assign _c_characterGenerator[3966] = 8'h00;
assign _c_characterGenerator[3967] = 8'h00;
assign _c_characterGenerator[3968] = 8'h00;
assign _c_characterGenerator[3969] = 8'h38;
assign _c_characterGenerator[3970] = 8'h6c;
assign _c_characterGenerator[3971] = 8'h6c;
assign _c_characterGenerator[3972] = 8'h38;
assign _c_characterGenerator[3973] = 8'h00;
assign _c_characterGenerator[3974] = 8'h00;
assign _c_characterGenerator[3975] = 8'h00;
assign _c_characterGenerator[3976] = 8'h00;
assign _c_characterGenerator[3977] = 8'h00;
assign _c_characterGenerator[3978] = 8'h00;
assign _c_characterGenerator[3979] = 8'h00;
assign _c_characterGenerator[3980] = 8'h00;
assign _c_characterGenerator[3981] = 8'h00;
assign _c_characterGenerator[3982] = 8'h00;
assign _c_characterGenerator[3983] = 8'h00;
assign _c_characterGenerator[3984] = 8'h00;
assign _c_characterGenerator[3985] = 8'h00;
assign _c_characterGenerator[3986] = 8'h00;
assign _c_characterGenerator[3987] = 8'h00;
assign _c_characterGenerator[3988] = 8'h00;
assign _c_characterGenerator[3989] = 8'h00;
assign _c_characterGenerator[3990] = 8'h00;
assign _c_characterGenerator[3991] = 8'h18;
assign _c_characterGenerator[3992] = 8'h18;
assign _c_characterGenerator[3993] = 8'h00;
assign _c_characterGenerator[3994] = 8'h00;
assign _c_characterGenerator[3995] = 8'h00;
assign _c_characterGenerator[3996] = 8'h00;
assign _c_characterGenerator[3997] = 8'h00;
assign _c_characterGenerator[3998] = 8'h00;
assign _c_characterGenerator[3999] = 8'h00;
assign _c_characterGenerator[4000] = 8'h00;
assign _c_characterGenerator[4001] = 8'h00;
assign _c_characterGenerator[4002] = 8'h00;
assign _c_characterGenerator[4003] = 8'h00;
assign _c_characterGenerator[4004] = 8'h00;
assign _c_characterGenerator[4005] = 8'h00;
assign _c_characterGenerator[4006] = 8'h00;
assign _c_characterGenerator[4007] = 8'h00;
assign _c_characterGenerator[4008] = 8'h18;
assign _c_characterGenerator[4009] = 8'h00;
assign _c_characterGenerator[4010] = 8'h00;
assign _c_characterGenerator[4011] = 8'h00;
assign _c_characterGenerator[4012] = 8'h00;
assign _c_characterGenerator[4013] = 8'h00;
assign _c_characterGenerator[4014] = 8'h00;
assign _c_characterGenerator[4015] = 8'h00;
assign _c_characterGenerator[4016] = 8'h00;
assign _c_characterGenerator[4017] = 8'h0f;
assign _c_characterGenerator[4018] = 8'h0c;
assign _c_characterGenerator[4019] = 8'h0c;
assign _c_characterGenerator[4020] = 8'h0c;
assign _c_characterGenerator[4021] = 8'h0c;
assign _c_characterGenerator[4022] = 8'h0c;
assign _c_characterGenerator[4023] = 8'hec;
assign _c_characterGenerator[4024] = 8'h6c;
assign _c_characterGenerator[4025] = 8'h6c;
assign _c_characterGenerator[4026] = 8'h3c;
assign _c_characterGenerator[4027] = 8'h1c;
assign _c_characterGenerator[4028] = 8'h00;
assign _c_characterGenerator[4029] = 8'h00;
assign _c_characterGenerator[4030] = 8'h00;
assign _c_characterGenerator[4031] = 8'h00;
assign _c_characterGenerator[4032] = 8'h00;
assign _c_characterGenerator[4033] = 8'hd8;
assign _c_characterGenerator[4034] = 8'h6c;
assign _c_characterGenerator[4035] = 8'h6c;
assign _c_characterGenerator[4036] = 8'h6c;
assign _c_characterGenerator[4037] = 8'h6c;
assign _c_characterGenerator[4038] = 8'h6c;
assign _c_characterGenerator[4039] = 8'h00;
assign _c_characterGenerator[4040] = 8'h00;
assign _c_characterGenerator[4041] = 8'h00;
assign _c_characterGenerator[4042] = 8'h00;
assign _c_characterGenerator[4043] = 8'h00;
assign _c_characterGenerator[4044] = 8'h00;
assign _c_characterGenerator[4045] = 8'h00;
assign _c_characterGenerator[4046] = 8'h00;
assign _c_characterGenerator[4047] = 8'h00;
assign _c_characterGenerator[4048] = 8'h00;
assign _c_characterGenerator[4049] = 8'h70;
assign _c_characterGenerator[4050] = 8'hd8;
assign _c_characterGenerator[4051] = 8'h30;
assign _c_characterGenerator[4052] = 8'h60;
assign _c_characterGenerator[4053] = 8'hc8;
assign _c_characterGenerator[4054] = 8'hf8;
assign _c_characterGenerator[4055] = 8'h00;
assign _c_characterGenerator[4056] = 8'h00;
assign _c_characterGenerator[4057] = 8'h00;
assign _c_characterGenerator[4058] = 8'h00;
assign _c_characterGenerator[4059] = 8'h00;
assign _c_characterGenerator[4060] = 8'h00;
assign _c_characterGenerator[4061] = 8'h00;
assign _c_characterGenerator[4062] = 8'h00;
assign _c_characterGenerator[4063] = 8'h00;
assign _c_characterGenerator[4064] = 8'h00;
assign _c_characterGenerator[4065] = 8'h00;
assign _c_characterGenerator[4066] = 8'h00;
assign _c_characterGenerator[4067] = 8'h00;
assign _c_characterGenerator[4068] = 8'h7c;
assign _c_characterGenerator[4069] = 8'h7c;
assign _c_characterGenerator[4070] = 8'h7c;
assign _c_characterGenerator[4071] = 8'h7c;
assign _c_characterGenerator[4072] = 8'h7c;
assign _c_characterGenerator[4073] = 8'h7c;
assign _c_characterGenerator[4074] = 8'h7c;
assign _c_characterGenerator[4075] = 8'h00;
assign _c_characterGenerator[4076] = 8'h00;
assign _c_characterGenerator[4077] = 8'h00;
assign _c_characterGenerator[4078] = 8'h00;
assign _c_characterGenerator[4079] = 8'h00;
assign _c_characterGenerator[4080] = 8'h00;
assign _c_characterGenerator[4081] = 8'h00;
assign _c_characterGenerator[4082] = 8'h00;
assign _c_characterGenerator[4083] = 8'h00;
assign _c_characterGenerator[4084] = 8'h00;
assign _c_characterGenerator[4085] = 8'h00;
assign _c_characterGenerator[4086] = 8'h00;
assign _c_characterGenerator[4087] = 8'h00;
assign _c_characterGenerator[4088] = 8'h00;
assign _c_characterGenerator[4089] = 8'h00;
assign _c_characterGenerator[4090] = 8'h00;
assign _c_characterGenerator[4091] = 8'h00;
assign _c_characterGenerator[4092] = 8'h00;
assign _c_characterGenerator[4093] = 8'h00;
assign _c_characterGenerator[4094] = 8'h00;
assign _c_characterGenerator[4095] = 8'h00;
wire  [7:0] _c_character_wdata0;
assign _c_character_wdata0 = 0;
wire  [7:0] _c_foreground_wdata0;
assign _c_foreground_wdata0 = 0;
wire  [7:0] _c_background_wdata0;
assign _c_background_wdata0 = 0;
wire  [7:0] _c_bitmap_wdata0;
assign _c_bitmap_wdata0 = 0;
wire  [5:0] _c_colourexpand3to6[7:0];
assign _c_colourexpand3to6[0] = 0;
assign _c_colourexpand3to6[1] = 9;
assign _c_colourexpand3to6[2] = 18;
assign _c_colourexpand3to6[3] = 27;
assign _c_colourexpand3to6[4] = 36;
assign _c_colourexpand3to6[5] = 45;
assign _c_colourexpand3to6[6] = 54;
assign _c_colourexpand3to6[7] = 63;
wire  [5:0] _c_colourexpand2to6[3:0];
assign _c_colourexpand2to6[0] = 0;
assign _c_colourexpand2to6[1] = 21;
assign _c_colourexpand2to6[2] = 42;
assign _c_colourexpand2to6[3] = 63;
wire  [7:0] _w_xcharacterpos;
wire  [11:0] _w_ycharacterpos;
wire  [7:0] _w_xincharacter;
wire  [7:0] _w_yincharacter;
wire  [0:0] _w_characterpixel;

reg  [0:0] _d_character_wenable0;
reg  [0:0] _q_character_wenable0;
reg  [11:0] _d_character_addr0;
reg  [11:0] _q_character_addr0;
reg  [0:0] _d_character_wenable1;
reg  [0:0] _q_character_wenable1;
reg  [7:0] _d_character_wdata1;
reg  [7:0] _q_character_wdata1;
reg  [11:0] _d_character_addr1;
reg  [11:0] _q_character_addr1;
reg  [0:0] _d_foreground_wenable0;
reg  [0:0] _q_foreground_wenable0;
reg  [11:0] _d_foreground_addr0;
reg  [11:0] _q_foreground_addr0;
reg  [0:0] _d_foreground_wenable1;
reg  [0:0] _q_foreground_wenable1;
reg  [7:0] _d_foreground_wdata1;
reg  [7:0] _q_foreground_wdata1;
reg  [11:0] _d_foreground_addr1;
reg  [11:0] _q_foreground_addr1;
reg  [0:0] _d_background_wenable0;
reg  [0:0] _q_background_wenable0;
reg  [11:0] _d_background_addr0;
reg  [11:0] _q_background_addr0;
reg  [0:0] _d_background_wenable1;
reg  [0:0] _q_background_wenable1;
reg  [7:0] _d_background_wdata1;
reg  [7:0] _q_background_wdata1;
reg  [11:0] _d_background_addr1;
reg  [11:0] _q_background_addr1;
reg  [0:0] _d_bitmap_wenable0;
reg  [0:0] _q_bitmap_wenable0;
reg  [18:0] _d_bitmap_addr0;
reg  [18:0] _q_bitmap_addr0;
reg  [0:0] _d_bitmap_wenable1;
reg  [0:0] _q_bitmap_wenable1;
reg  [7:0] _d_bitmap_wdata1;
reg  [7:0] _q_bitmap_wdata1;
reg  [18:0] _d_bitmap_addr1;
reg  [18:0] _q_bitmap_addr1;
reg  [5:0] _d_pix_red,_q_pix_red;
reg  [5:0] _d_pix_green,_q_pix_green;
reg  [5:0] _d_pix_blue,_q_pix_blue;
reg  [1:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_character_wenable0 <= 0;
_q_character_addr0 <= 0;
_q_character_wenable1 <= 0;
_q_character_wdata1 <= 0;
_q_character_addr1 <= 0;
_q_foreground_wenable0 <= 0;
_q_foreground_addr0 <= 0;
_q_foreground_wenable1 <= 0;
_q_foreground_wdata1 <= 0;
_q_foreground_addr1 <= 0;
_q_background_wenable0 <= 0;
_q_background_addr0 <= 0;
_q_background_wenable1 <= 0;
_q_background_wdata1 <= 0;
_q_background_addr1 <= 0;
_q_bitmap_wenable0 <= 0;
_q_bitmap_addr0 <= 0;
_q_bitmap_wenable1 <= 0;
_q_bitmap_wdata1 <= 0;
_q_bitmap_addr1 <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_character_wenable0 <= _d_character_wenable0;
_q_character_addr0 <= _d_character_addr0;
_q_character_wenable1 <= _d_character_wenable1;
_q_character_wdata1 <= _d_character_wdata1;
_q_character_addr1 <= _d_character_addr1;
_q_foreground_wenable0 <= _d_foreground_wenable0;
_q_foreground_addr0 <= _d_foreground_addr0;
_q_foreground_wenable1 <= _d_foreground_wenable1;
_q_foreground_wdata1 <= _d_foreground_wdata1;
_q_foreground_addr1 <= _d_foreground_addr1;
_q_background_wenable0 <= _d_background_wenable0;
_q_background_addr0 <= _d_background_addr0;
_q_background_wenable1 <= _d_background_wenable1;
_q_background_wdata1 <= _d_background_wdata1;
_q_background_addr1 <= _d_background_addr1;
_q_bitmap_wenable0 <= _d_bitmap_wenable0;
_q_bitmap_addr0 <= _d_bitmap_addr0;
_q_bitmap_wenable1 <= _d_bitmap_wenable1;
_q_bitmap_wdata1 <= _d_bitmap_wdata1;
_q_bitmap_addr1 <= _d_bitmap_addr1;
_q_index <= _d_index;
  end
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
end


M_multiplex_display_mem_character __mem__character(
.clock0(clock),
.clock1(clock),
.in_character_wenable0(_d_character_wenable0),
.in_character_wdata0(_c_character_wdata0),
.in_character_addr0(_d_character_addr0),
.in_character_wenable1(_d_character_wenable1),
.in_character_wdata1(_d_character_wdata1),
.in_character_addr1(_d_character_addr1),
.out_character_rdata0(_w_mem_character_rdata0),
.out_character_rdata1(_w_mem_character_rdata1)
);
M_multiplex_display_mem_foreground __mem__foreground(
.clock0(clock),
.clock1(clock),
.in_foreground_wenable0(_d_foreground_wenable0),
.in_foreground_wdata0(_c_foreground_wdata0),
.in_foreground_addr0(_d_foreground_addr0),
.in_foreground_wenable1(_d_foreground_wenable1),
.in_foreground_wdata1(_d_foreground_wdata1),
.in_foreground_addr1(_d_foreground_addr1),
.out_foreground_rdata0(_w_mem_foreground_rdata0),
.out_foreground_rdata1(_w_mem_foreground_rdata1)
);
M_multiplex_display_mem_background __mem__background(
.clock0(clock),
.clock1(clock),
.in_background_wenable0(_d_background_wenable0),
.in_background_wdata0(_c_background_wdata0),
.in_background_addr0(_d_background_addr0),
.in_background_wenable1(_d_background_wenable1),
.in_background_wdata1(_d_background_wdata1),
.in_background_addr1(_d_background_addr1),
.out_background_rdata0(_w_mem_background_rdata0),
.out_background_rdata1(_w_mem_background_rdata1)
);
M_multiplex_display_mem_bitmap __mem__bitmap(
.clock0(clock),
.clock1(clock),
.in_bitmap_wenable0(_d_bitmap_wenable0),
.in_bitmap_wdata0(_c_bitmap_wdata0),
.in_bitmap_addr0(_d_bitmap_addr0),
.in_bitmap_wenable1(_d_bitmap_wenable1),
.in_bitmap_wdata1(_d_bitmap_wdata1),
.in_bitmap_addr1(_d_bitmap_addr1),
.out_bitmap_rdata0(_w_mem_bitmap_rdata0),
.out_bitmap_rdata1(_w_mem_bitmap_rdata1)
);

assign _w_characterpixel = ((_c_characterGenerator[_w_mem_character_rdata0*16+_w_yincharacter]<<_w_xincharacter)>>7)&1;
assign _w_yincharacter = in_pix_y&15;
assign _w_ycharacterpos = ((in_pix_y)>>4)*80;
assign _w_xincharacter = in_pix_x&7;
assign _w_xcharacterpos = (in_pix_x+1)>>3;

always @* begin
_d_character_wenable0 = _q_character_wenable0;
_d_character_addr0 = _q_character_addr0;
_d_character_wenable1 = _q_character_wenable1;
_d_character_wdata1 = _q_character_wdata1;
_d_character_addr1 = _q_character_addr1;
_d_foreground_wenable0 = _q_foreground_wenable0;
_d_foreground_addr0 = _q_foreground_addr0;
_d_foreground_wenable1 = _q_foreground_wenable1;
_d_foreground_wdata1 = _q_foreground_wdata1;
_d_foreground_addr1 = _q_foreground_addr1;
_d_background_wenable0 = _q_background_wenable0;
_d_background_addr0 = _q_background_addr0;
_d_background_wenable1 = _q_background_wenable1;
_d_background_wdata1 = _q_background_wdata1;
_d_background_addr1 = _q_background_addr1;
_d_bitmap_wenable0 = _q_bitmap_wenable0;
_d_bitmap_addr0 = _q_bitmap_addr0;
_d_bitmap_wenable1 = _q_bitmap_wenable1;
_d_bitmap_wdata1 = _q_bitmap_wdata1;
_d_bitmap_addr1 = _q_bitmap_addr1;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_index = _q_index;
// _always_pre
_d_pix_red = 0;
_d_pix_green = 0;
_d_pix_blue = 0;
_d_character_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_character_wenable0 = 0;
_d_foreground_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_foreground_wenable0 = 0;
_d_background_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_background_wenable0 = 0;
_d_bitmap_addr0 = in_pix_x+in_pix_y*640;
_d_bitmap_wenable0 = 0;
_d_bitmap_addr1 = in_gpu_x+in_gpu_y*640;
_d_bitmap_wenable1 = 0;
_d_character_addr1 = in_tpu_x+in_tpu_y*80;
_d_character_wenable1 = 0;
_d_background_addr1 = in_tpu_x+in_tpu_y*80;
_d_background_wenable1 = 0;
_d_foreground_addr1 = in_tpu_x+in_tpu_y*80;
_d_foreground_wenable1 = 0;
_d_index = 3;
case (_q_index)
0: begin
// _top
// var inits
_d_character_wenable0 = 0;
_d_character_addr0 = 0;
_d_character_wenable1 = 0;
_d_character_wdata1 = 0;
_d_character_addr1 = 0;
_d_foreground_wenable0 = 0;
_d_foreground_addr0 = 0;
_d_foreground_wenable1 = 0;
_d_foreground_wdata1 = 0;
_d_foreground_addr1 = 0;
_d_background_wenable0 = 0;
_d_background_addr0 = 0;
_d_background_wenable1 = 0;
_d_background_wdata1 = 0;
_d_background_addr1 = 0;
_d_bitmap_wenable0 = 0;
_d_bitmap_addr0 = 0;
_d_bitmap_wenable1 = 0;
_d_bitmap_wdata1 = 0;
_d_bitmap_addr1 = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_gpu_write) begin
// __block_5
// __block_7
_d_bitmap_wdata1 = in_gpu_dotset;
_d_bitmap_wenable1 = 1;
// __block_8
end else begin
// __block_6
end
// __block_9
  case (in_tpu_write)
  1: begin
// __block_11_case
// __block_12
_d_character_wdata1 = in_tpu_set;
_d_character_wenable1 = 1;
// __block_13
  end
  2: begin
// __block_14_case
// __block_15
_d_background_wdata1 = in_tpu_set;
_d_background_wenable1 = 1;
// __block_16
  end
  3: begin
// __block_17_case
// __block_18
_d_foreground_wdata1 = in_tpu_set;
_d_foreground_wenable1 = 1;
// __block_19
  end
  default: begin
// __block_20_case
// __block_21
// __block_22
  end
endcase
// __block_10
if (in_pix_vblank==0) begin
// __block_23
// __block_25
if (in_pix_active) begin
// __block_26
// __block_28
  case (_w_mem_character_rdata0)
  0: begin
// __block_30_case
// __block_31
_d_pix_red = _c_colourexpand3to6[(_w_mem_bitmap_rdata0&8'he0)>>5];
_d_pix_green = _c_colourexpand3to6[(_w_mem_bitmap_rdata0&8'h1c)>>2];
_d_pix_blue = _c_colourexpand2to6[(_w_mem_bitmap_rdata0&8'h3)];
// __block_32
  end
  default: begin
// __block_33_case
// __block_34
  case (_w_characterpixel)
  0: begin
// __block_36_case
// __block_37
_d_pix_red = _c_colourexpand3to6[(_w_mem_background_rdata0&8'he0)>>5];
_d_pix_green = _c_colourexpand3to6[(_w_mem_background_rdata0&8'h1c)>>2];
_d_pix_blue = _c_colourexpand2to6[(_w_mem_background_rdata0&8'h3)];
// __block_38
  end
  1: begin
// __block_39_case
// __block_40
_d_pix_red = _c_colourexpand3to6[(_w_mem_foreground_rdata0&8'he0)>>5];
_d_pix_green = _c_colourexpand3to6[(_w_mem_foreground_rdata0&8'h1c)>>2];
_d_pix_blue = _c_colourexpand2to6[(_w_mem_foreground_rdata0&8'h3)];
// __block_41
  end
endcase
// __block_35
// __block_42
  end
endcase
// __block_29
// __block_43
end else begin
// __block_27
end
// __block_44
// __block_45
end else begin
// __block_24
end
// __block_46
// __block_47
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of multiplex_display
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_main_mem_dstack(
input                  [0:0] in_dstack_wenable,
input       [15:0]    in_dstack_wdata,
input                  [7:0]    in_dstack_addr,
output reg  [15:0]    out_dstack_rdata,
input                                      clock
);
reg  [15:0] buffer[255:0];
always @(posedge clock) begin
  if (in_dstack_wenable) begin
    buffer[in_dstack_addr] <= in_dstack_wdata;
  end
  out_dstack_rdata <= buffer[in_dstack_addr];
end

endmodule

module M_main_mem_rstack(
input                  [0:0] in_rstack_wenable,
input       [15:0]    in_rstack_wdata,
input                  [7:0]    in_rstack_addr,
output reg  [15:0]    out_rstack_rdata,
input                                      clock
);
reg  [15:0] buffer[255:0];
always @(posedge clock) begin
  if (in_rstack_wenable) begin
    buffer[in_rstack_addr] <= in_rstack_wdata;
  end
  out_rstack_rdata <= buffer[in_rstack_addr];
end

endmodule

module M_main_mem_rom(
input                  [11:0] in_rom_addr,
output reg  [15:0] out_rom_rdata,
input                                   clock
);
reg  [15:0] buffer[3652:0];
always @(posedge clock) begin
   out_rom_rdata <= buffer[in_rom_addr];
end
initial begin
 buffer[0] = 16'h0E2D;
 buffer[1] = 16'h0010;
 buffer[2] = 16'h0000;
 buffer[3] = 16'h0000;
 buffer[4] = 16'h0000;
 buffer[5] = 16'h7F00;
 buffer[6] = 16'h10AE;
 buffer[7] = 16'h118C;
 buffer[8] = 16'h0000;
 buffer[9] = 16'h0000;
 buffer[10] = 16'h0000;
 buffer[11] = 16'h0000;
 buffer[12] = 16'h0000;
 buffer[13] = 16'h0000;
 buffer[14] = 16'h0000;
 buffer[15] = 16'h0000;
 buffer[16] = 16'h0000;
 buffer[17] = 16'h0000;
 buffer[18] = 16'h0000;
 buffer[19] = 16'h0000;
 buffer[20] = 16'h0000;
 buffer[21] = 16'h0000;
 buffer[22] = 16'h0000;
 buffer[23] = 16'h1C8A;
 buffer[24] = 16'h1C54;
 buffer[25] = 16'h0952;
 buffer[26] = 16'h0964;
 buffer[27] = 16'h1C20;
 buffer[28] = 16'h0E6A;
 buffer[29] = 16'h0F56;
 buffer[30] = 16'h1662;
 buffer[31] = 16'h16E4;
 buffer[32] = 16'h170C;
 buffer[33] = 16'h1778;
 buffer[34] = 16'h0000;
 buffer[35] = 16'h0000;
 buffer[36] = 16'h0000;
 buffer[37] = 16'h0000;
 buffer[38] = 16'h0000;
 buffer[39] = 16'h0000;
 buffer[40] = 16'h0000;
 buffer[41] = 16'h0000;
 buffer[42] = 16'h0000;
 buffer[43] = 16'h0000;
 buffer[44] = 16'h0000;
 buffer[45] = 16'h0000;
 buffer[46] = 16'h0000;
 buffer[47] = 16'h0000;
 buffer[48] = 16'h0000;
 buffer[49] = 16'h0000;
 buffer[50] = 16'h0000;
 buffer[51] = 16'h0000;
 buffer[52] = 16'h0000;
 buffer[53] = 16'h0000;
 buffer[54] = 16'h0000;
 buffer[55] = 16'h0000;
 buffer[56] = 16'h0000;
 buffer[57] = 16'h0000;
 buffer[58] = 16'h0000;
 buffer[59] = 16'h0000;
 buffer[60] = 16'h0000;
 buffer[61] = 16'h0000;
 buffer[62] = 16'h0000;
 buffer[63] = 16'h0000;
 buffer[64] = 16'h6003;
 buffer[65] = 16'h6003;
 buffer[66] = 16'h6003;
 buffer[67] = 16'h6003;
 buffer[68] = 16'h6003;
 buffer[69] = 16'h6003;
 buffer[70] = 16'h6003;
 buffer[71] = 16'h6003;
 buffer[72] = 16'h6003;
 buffer[73] = 16'h6003;
 buffer[74] = 16'h6003;
 buffer[75] = 16'h6003;
 buffer[76] = 16'h6003;
 buffer[77] = 16'h6003;
 buffer[78] = 16'h6003;
 buffer[79] = 16'h710C;
 buffer[80] = 16'h6001;
 buffer[81] = 16'h6001;
 buffer[82] = 16'h6001;
 buffer[83] = 16'h6001;
 buffer[84] = 16'h6001;
 buffer[85] = 16'h6001;
 buffer[86] = 16'h6001;
 buffer[87] = 16'h6001;
 buffer[88] = 16'h6001;
 buffer[89] = 16'h6001;
 buffer[90] = 16'h6001;
 buffer[91] = 16'h6001;
 buffer[92] = 16'h6001;
 buffer[93] = 16'h6001;
 buffer[94] = 16'h6001;
 buffer[95] = 16'h700C;
 buffer[96] = 16'h6100;
 buffer[97] = 16'h700C;
 buffer[98] = 16'h404E;
 buffer[99] = 16'h005E;
 buffer[100] = 16'h404D;
 buffer[101] = 16'h005D;
 buffer[102] = 16'h404C;
 buffer[103] = 16'h005C;
 buffer[104] = 16'h404B;
 buffer[105] = 16'h005B;
 buffer[106] = 16'h404A;
 buffer[107] = 16'h005A;
 buffer[108] = 16'h4049;
 buffer[109] = 16'h0059;
 buffer[110] = 16'h4048;
 buffer[111] = 16'h0058;
 buffer[112] = 16'h4047;
 buffer[113] = 16'h0057;
 buffer[114] = 16'h4046;
 buffer[115] = 16'h0056;
 buffer[116] = 16'h4045;
 buffer[117] = 16'h0055;
 buffer[118] = 16'h4044;
 buffer[119] = 16'h0054;
 buffer[120] = 16'h4043;
 buffer[121] = 16'h0053;
 buffer[122] = 16'h4042;
 buffer[123] = 16'h0052;
 buffer[124] = 16'h4041;
 buffer[125] = 16'h0051;
 buffer[126] = 16'h4040;
 buffer[127] = 16'h0050;
 buffer[128] = 16'h700C;
 buffer[129] = 16'h0000;
 buffer[130] = 16'h0000;
 buffer[131] = 16'h0000;
 buffer[132] = 16'h0000;
 buffer[133] = 16'h0000;
 buffer[134] = 16'h0000;
 buffer[135] = 16'h0000;
 buffer[136] = 16'h0000;
 buffer[137] = 16'h0000;
 buffer[138] = 16'h0000;
 buffer[139] = 16'h0000;
 buffer[140] = 16'h0000;
 buffer[141] = 16'h0000;
 buffer[142] = 16'h0000;
 buffer[143] = 16'h0000;
 buffer[144] = 16'h0000;
 buffer[145] = 16'h0000;
 buffer[146] = 16'h0000;
 buffer[147] = 16'h0000;
 buffer[148] = 16'h0000;
 buffer[149] = 16'h0000;
 buffer[150] = 16'h0000;
 buffer[151] = 16'h0000;
 buffer[152] = 16'h0000;
 buffer[153] = 16'h0000;
 buffer[154] = 16'h0000;
 buffer[155] = 16'h0000;
 buffer[156] = 16'h0000;
 buffer[157] = 16'h0000;
 buffer[158] = 16'h0000;
 buffer[159] = 16'h0000;
 buffer[160] = 16'h0000;
 buffer[161] = 16'h0000;
 buffer[162] = 16'h0000;
 buffer[163] = 16'h0000;
 buffer[164] = 16'h0000;
 buffer[165] = 16'h0000;
 buffer[166] = 16'h0000;
 buffer[167] = 16'h0000;
 buffer[168] = 16'h0000;
 buffer[169] = 16'h0000;
 buffer[170] = 16'h0000;
 buffer[171] = 16'h0000;
 buffer[172] = 16'h0000;
 buffer[173] = 16'h0000;
 buffer[174] = 16'h0000;
 buffer[175] = 16'h0000;
 buffer[176] = 16'h0000;
 buffer[177] = 16'h0000;
 buffer[178] = 16'h0000;
 buffer[179] = 16'h0000;
 buffer[180] = 16'h0000;
 buffer[181] = 16'h0000;
 buffer[182] = 16'h0000;
 buffer[183] = 16'h0000;
 buffer[184] = 16'h0000;
 buffer[185] = 16'h0000;
 buffer[186] = 16'h0000;
 buffer[187] = 16'h0000;
 buffer[188] = 16'h0000;
 buffer[189] = 16'h0000;
 buffer[190] = 16'h0000;
 buffer[191] = 16'h0000;
 buffer[192] = 16'h0000;
 buffer[193] = 16'h6E04;
 buffer[194] = 16'h6F6F;
 buffer[195] = 16'h0070;
 buffer[196] = 16'h700C;
 buffer[197] = 16'h0182;
 buffer[198] = 16'h2B01;
 buffer[199] = 16'h720F;
 buffer[200] = 16'h018C;
 buffer[201] = 16'h7803;
 buffer[202] = 16'h726F;
 buffer[203] = 16'h750F;
 buffer[204] = 16'h0192;
 buffer[205] = 16'h6103;
 buffer[206] = 16'h646E;
 buffer[207] = 16'h730F;
 buffer[208] = 16'h019A;
 buffer[209] = 16'h6F02;
 buffer[210] = 16'h0072;
 buffer[211] = 16'h740F;
 buffer[212] = 16'h01A2;
 buffer[213] = 16'h6906;
 buffer[214] = 16'h766E;
 buffer[215] = 16'h7265;
 buffer[216] = 16'h0074;
 buffer[217] = 16'h760C;
 buffer[218] = 16'h01AA;
 buffer[219] = 16'h3D01;
 buffer[220] = 16'h770F;
 buffer[221] = 16'h01B6;
 buffer[222] = 16'h3C01;
 buffer[223] = 16'h780F;
 buffer[224] = 16'h01BC;
 buffer[225] = 16'h7502;
 buffer[226] = 16'h003C;
 buffer[227] = 16'h7F0F;
 buffer[228] = 16'h01C2;
 buffer[229] = 16'h7304;
 buffer[230] = 16'h6177;
 buffer[231] = 16'h0070;
 buffer[232] = 16'h718C;
 buffer[233] = 16'h01CA;
 buffer[234] = 16'h7502;
 buffer[235] = 16'h003E;
 buffer[236] = 16'h771F;
 buffer[237] = 16'h01D4;
 buffer[238] = 16'h6403;
 buffer[239] = 16'h7075;
 buffer[240] = 16'h708D;
 buffer[241] = 16'h01DC;
 buffer[242] = 16'h6404;
 buffer[243] = 16'h6F72;
 buffer[244] = 16'h0070;
 buffer[245] = 16'h710F;
 buffer[246] = 16'h01E4;
 buffer[247] = 16'h6F04;
 buffer[248] = 16'h6576;
 buffer[249] = 16'h0072;
 buffer[250] = 16'h718D;
 buffer[251] = 16'h01EE;
 buffer[252] = 16'h6E03;
 buffer[253] = 16'h7069;
 buffer[254] = 16'h700F;
 buffer[255] = 16'h01F8;
 buffer[256] = 16'h6C06;
 buffer[257] = 16'h6873;
 buffer[258] = 16'h6669;
 buffer[259] = 16'h0074;
 buffer[260] = 16'h7D0F;
 buffer[261] = 16'h0200;
 buffer[262] = 16'h7206;
 buffer[263] = 16'h6873;
 buffer[264] = 16'h6669;
 buffer[265] = 16'h0074;
 buffer[266] = 16'h790F;
 buffer[267] = 16'h020C;
 buffer[268] = 16'h3102;
 buffer[269] = 16'h002D;
 buffer[270] = 16'h7A0C;
 buffer[271] = 16'h0218;
 buffer[272] = 16'h3E42;
 buffer[273] = 16'h0072;
 buffer[274] = 16'h6B8D;
 buffer[275] = 16'h6180;
 buffer[276] = 16'h6147;
 buffer[277] = 16'h6147;
 buffer[278] = 16'h700C;
 buffer[279] = 16'h0220;
 buffer[280] = 16'h7242;
 buffer[281] = 16'h003E;
 buffer[282] = 16'h6B8D;
 buffer[283] = 16'h6B8D;
 buffer[284] = 16'h6180;
 buffer[285] = 16'h6147;
 buffer[286] = 16'h700C;
 buffer[287] = 16'h0230;
 buffer[288] = 16'h7242;
 buffer[289] = 16'h0040;
 buffer[290] = 16'h6B8D;
 buffer[291] = 16'h6B8D;
 buffer[292] = 16'h6081;
 buffer[293] = 16'h6147;
 buffer[294] = 16'h6180;
 buffer[295] = 16'h6147;
 buffer[296] = 16'h700C;
 buffer[297] = 16'h0240;
 buffer[298] = 16'h4001;
 buffer[299] = 16'h7C0C;
 buffer[300] = 16'h0254;
 buffer[301] = 16'h2101;
 buffer[302] = 16'h6023;
 buffer[303] = 16'h710F;
 buffer[304] = 16'h025A;
 buffer[305] = 16'h3C02;
 buffer[306] = 16'h003E;
 buffer[307] = 16'h721F;
 buffer[308] = 16'h0262;
 buffer[309] = 16'h3002;
 buffer[310] = 16'h003C;
 buffer[311] = 16'h781C;
 buffer[312] = 16'h026A;
 buffer[313] = 16'h3002;
 buffer[314] = 16'h003D;
 buffer[315] = 16'h701C;
 buffer[316] = 16'h0272;
 buffer[317] = 16'h3003;
 buffer[318] = 16'h3E3C;
 buffer[319] = 16'h711C;
 buffer[320] = 16'h027A;
 buffer[321] = 16'h3E01;
 buffer[322] = 16'h761F;
 buffer[323] = 16'h0282;
 buffer[324] = 16'h3002;
 buffer[325] = 16'h003E;
 buffer[326] = 16'h791C;
 buffer[327] = 16'h0288;
 buffer[328] = 16'h3E02;
 buffer[329] = 16'h003D;
 buffer[330] = 16'h7F1F;
 buffer[331] = 16'h0290;
 buffer[332] = 16'h7404;
 buffer[333] = 16'h6375;
 buffer[334] = 16'h006B;
 buffer[335] = 16'h6180;
 buffer[336] = 16'h718D;
 buffer[337] = 16'h0298;
 buffer[338] = 16'h2D04;
 buffer[339] = 16'h6F72;
 buffer[340] = 16'h0074;
 buffer[341] = 16'h6180;
 buffer[342] = 16'h6147;
 buffer[343] = 16'h6180;
 buffer[344] = 16'h6B8D;
 buffer[345] = 16'h700C;
 buffer[346] = 16'h02A4;
 buffer[347] = 16'h3202;
 buffer[348] = 16'h002F;
 buffer[349] = 16'h8001;
 buffer[350] = 16'h790F;
 buffer[351] = 16'h02B6;
 buffer[352] = 16'h3202;
 buffer[353] = 16'h002A;
 buffer[354] = 16'h741C;
 buffer[355] = 16'h02C0;
 buffer[356] = 16'h3102;
 buffer[357] = 16'h002B;
 buffer[358] = 16'h731C;
 buffer[359] = 16'h02C8;
 buffer[360] = 16'h7303;
 buffer[361] = 16'h4070;
 buffer[362] = 16'h6E81;
 buffer[363] = 16'h80FF;
 buffer[364] = 16'h730F;
 buffer[365] = 16'h02D0;
 buffer[366] = 16'h6507;
 buffer[367] = 16'h6578;
 buffer[368] = 16'h7563;
 buffer[369] = 16'h6574;
 buffer[370] = 16'h6147;
 buffer[371] = 16'h700C;
 buffer[372] = 16'h02DC;
 buffer[373] = 16'h6203;
 buffer[374] = 16'h6579;
 buffer[375] = 16'h8FFD;
 buffer[376] = 16'h6600;
 buffer[377] = 16'h6023;
 buffer[378] = 16'h710F;
 buffer[379] = 16'h02EA;
 buffer[380] = 16'h6302;
 buffer[381] = 16'h0040;
 buffer[382] = 16'h6081;
 buffer[383] = 16'h6C00;
 buffer[384] = 16'h6180;
 buffer[385] = 16'h8001;
 buffer[386] = 16'h6303;
 buffer[387] = 16'h2187;
 buffer[388] = 16'h8008;
 buffer[389] = 16'h6903;
 buffer[390] = 16'h0189;
 buffer[391] = 16'h80FF;
 buffer[392] = 16'h730F;
 buffer[393] = 16'h700C;
 buffer[394] = 16'h02F8;
 buffer[395] = 16'h6302;
 buffer[396] = 16'h0021;
 buffer[397] = 16'h6180;
 buffer[398] = 16'h80FF;
 buffer[399] = 16'h6303;
 buffer[400] = 16'h6081;
 buffer[401] = 16'h8008;
 buffer[402] = 16'h6D03;
 buffer[403] = 16'h6403;
 buffer[404] = 16'h6180;
 buffer[405] = 16'h414F;
 buffer[406] = 16'h6081;
 buffer[407] = 16'h6C00;
 buffer[408] = 16'h6180;
 buffer[409] = 16'h8001;
 buffer[410] = 16'h6303;
 buffer[411] = 16'h8000;
 buffer[412] = 16'h6703;
 buffer[413] = 16'h80FF;
 buffer[414] = 16'h6503;
 buffer[415] = 16'h6147;
 buffer[416] = 16'h6181;
 buffer[417] = 16'h6503;
 buffer[418] = 16'h6B8D;
 buffer[419] = 16'h6303;
 buffer[420] = 16'h6503;
 buffer[421] = 16'h6180;
 buffer[422] = 16'h6023;
 buffer[423] = 16'h710F;
 buffer[424] = 16'h0316;
 buffer[425] = 16'h7503;
 buffer[426] = 16'h2B6D;
 buffer[427] = 16'h6181;
 buffer[428] = 16'h6181;
 buffer[429] = 16'h6203;
 buffer[430] = 16'h6147;
 buffer[431] = 16'h6B81;
 buffer[432] = 16'h8000;
 buffer[433] = 16'h6F13;
 buffer[434] = 16'h6147;
 buffer[435] = 16'h6181;
 buffer[436] = 16'h6181;
 buffer[437] = 16'h6303;
 buffer[438] = 16'h6810;
 buffer[439] = 16'h6B8D;
 buffer[440] = 16'h6403;
 buffer[441] = 16'h6147;
 buffer[442] = 16'h6403;
 buffer[443] = 16'h6810;
 buffer[444] = 16'h6B8D;
 buffer[445] = 16'h6303;
 buffer[446] = 16'h6600;
 buffer[447] = 16'h6310;
 buffer[448] = 16'h6B8D;
 buffer[449] = 16'h718C;
 buffer[450] = 16'h0352;
 buffer[451] = 16'h6445;
 buffer[452] = 16'h766F;
 buffer[453] = 16'h7261;
 buffer[454] = 16'h6B8D;
 buffer[455] = 16'h700C;
 buffer[456] = 16'h0386;
 buffer[457] = 16'h7502;
 buffer[458] = 16'h0070;
 buffer[459] = 16'h41C6;
 buffer[460] = 16'h7E8C;
 buffer[461] = 16'h0392;
 buffer[462] = 16'h6446;
 buffer[463] = 16'h756F;
 buffer[464] = 16'h6573;
 buffer[465] = 16'h0072;
 buffer[466] = 16'h41CB;
 buffer[467] = 16'h6C00;
 buffer[468] = 16'h6B8D;
 buffer[469] = 16'h6C00;
 buffer[470] = 16'h720F;
 buffer[471] = 16'h039C;
 buffer[472] = 16'h6204;
 buffer[473] = 16'h7361;
 buffer[474] = 16'h0065;
 buffer[475] = 16'hFE80;
 buffer[476] = 16'h700C;
 buffer[477] = 16'h03B0;
 buffer[478] = 16'h7404;
 buffer[479] = 16'h6D65;
 buffer[480] = 16'h0070;
 buffer[481] = 16'hFE82;
 buffer[482] = 16'h700C;
 buffer[483] = 16'h03BC;
 buffer[484] = 16'h3E03;
 buffer[485] = 16'h6E69;
 buffer[486] = 16'hFE84;
 buffer[487] = 16'h700C;
 buffer[488] = 16'h03C8;
 buffer[489] = 16'h2304;
 buffer[490] = 16'h6974;
 buffer[491] = 16'h0062;
 buffer[492] = 16'hFE86;
 buffer[493] = 16'h700C;
 buffer[494] = 16'h03D2;
 buffer[495] = 16'h7403;
 buffer[496] = 16'h6269;
 buffer[497] = 16'hFE88;
 buffer[498] = 16'h700C;
 buffer[499] = 16'h03DE;
 buffer[500] = 16'h2705;
 buffer[501] = 16'h7665;
 buffer[502] = 16'h6C61;
 buffer[503] = 16'hFE8A;
 buffer[504] = 16'h700C;
 buffer[505] = 16'h03E8;
 buffer[506] = 16'h2706;
 buffer[507] = 16'h6261;
 buffer[508] = 16'h726F;
 buffer[509] = 16'h0074;
 buffer[510] = 16'hFE8C;
 buffer[511] = 16'h700C;
 buffer[512] = 16'h03F4;
 buffer[513] = 16'h6803;
 buffer[514] = 16'h646C;
 buffer[515] = 16'hFE8E;
 buffer[516] = 16'h700C;
 buffer[517] = 16'h0402;
 buffer[518] = 16'h6307;
 buffer[519] = 16'h6E6F;
 buffer[520] = 16'h6574;
 buffer[521] = 16'h7478;
 buffer[522] = 16'hFE90;
 buffer[523] = 16'h700C;
 buffer[524] = 16'h040C;
 buffer[525] = 16'h660E;
 buffer[526] = 16'h726F;
 buffer[527] = 16'h6874;
 buffer[528] = 16'h772D;
 buffer[529] = 16'h726F;
 buffer[530] = 16'h6C64;
 buffer[531] = 16'h7369;
 buffer[532] = 16'h0074;
 buffer[533] = 16'hFEA2;
 buffer[534] = 16'h700C;
 buffer[535] = 16'h041A;
 buffer[536] = 16'h6307;
 buffer[537] = 16'h7275;
 buffer[538] = 16'h6572;
 buffer[539] = 16'h746E;
 buffer[540] = 16'hFEA8;
 buffer[541] = 16'h700C;
 buffer[542] = 16'h0430;
 buffer[543] = 16'h6402;
 buffer[544] = 16'h0070;
 buffer[545] = 16'hFEAC;
 buffer[546] = 16'h700C;
 buffer[547] = 16'h043E;
 buffer[548] = 16'h6C04;
 buffer[549] = 16'h7361;
 buffer[550] = 16'h0074;
 buffer[551] = 16'hFEAE;
 buffer[552] = 16'h700C;
 buffer[553] = 16'h0448;
 buffer[554] = 16'h2705;
 buffer[555] = 16'h6B3F;
 buffer[556] = 16'h7965;
 buffer[557] = 16'hFEB0;
 buffer[558] = 16'h700C;
 buffer[559] = 16'h0454;
 buffer[560] = 16'h2705;
 buffer[561] = 16'h6D65;
 buffer[562] = 16'h7469;
 buffer[563] = 16'hFEB2;
 buffer[564] = 16'h700C;
 buffer[565] = 16'h0460;
 buffer[566] = 16'h2705;
 buffer[567] = 16'h6F62;
 buffer[568] = 16'h746F;
 buffer[569] = 16'hFEB4;
 buffer[570] = 16'h700C;
 buffer[571] = 16'h046C;
 buffer[572] = 16'h2702;
 buffer[573] = 16'h005C;
 buffer[574] = 16'hFEB6;
 buffer[575] = 16'h700C;
 buffer[576] = 16'h0478;
 buffer[577] = 16'h2706;
 buffer[578] = 16'h616E;
 buffer[579] = 16'h656D;
 buffer[580] = 16'h003F;
 buffer[581] = 16'hFEB8;
 buffer[582] = 16'h700C;
 buffer[583] = 16'h0482;
 buffer[584] = 16'h2704;
 buffer[585] = 16'h2C24;
 buffer[586] = 16'h006E;
 buffer[587] = 16'hFEBA;
 buffer[588] = 16'h700C;
 buffer[589] = 16'h0490;
 buffer[590] = 16'h2706;
 buffer[591] = 16'h766F;
 buffer[592] = 16'h7265;
 buffer[593] = 16'h0074;
 buffer[594] = 16'hFEBC;
 buffer[595] = 16'h700C;
 buffer[596] = 16'h049C;
 buffer[597] = 16'h2702;
 buffer[598] = 16'h003B;
 buffer[599] = 16'hFEBE;
 buffer[600] = 16'h700C;
 buffer[601] = 16'h04AA;
 buffer[602] = 16'h2707;
 buffer[603] = 16'h7263;
 buffer[604] = 16'h6165;
 buffer[605] = 16'h6574;
 buffer[606] = 16'hFEC0;
 buffer[607] = 16'h700C;
 buffer[608] = 16'h04B4;
 buffer[609] = 16'h3F04;
 buffer[610] = 16'h7564;
 buffer[611] = 16'h0070;
 buffer[612] = 16'h6081;
 buffer[613] = 16'h2267;
 buffer[614] = 16'h708D;
 buffer[615] = 16'h700C;
 buffer[616] = 16'h04C2;
 buffer[617] = 16'h7203;
 buffer[618] = 16'h746F;
 buffer[619] = 16'h6147;
 buffer[620] = 16'h6180;
 buffer[621] = 16'h6B8D;
 buffer[622] = 16'h718C;
 buffer[623] = 16'h04D2;
 buffer[624] = 16'h3205;
 buffer[625] = 16'h7264;
 buffer[626] = 16'h706F;
 buffer[627] = 16'h6103;
 buffer[628] = 16'h710F;
 buffer[629] = 16'h04E0;
 buffer[630] = 16'h3204;
 buffer[631] = 16'h7564;
 buffer[632] = 16'h0070;
 buffer[633] = 16'h6181;
 buffer[634] = 16'h718D;
 buffer[635] = 16'h04EC;
 buffer[636] = 16'h6E06;
 buffer[637] = 16'h6765;
 buffer[638] = 16'h7461;
 buffer[639] = 16'h0065;
 buffer[640] = 16'h7D1C;
 buffer[641] = 16'h04F8;
 buffer[642] = 16'h6407;
 buffer[643] = 16'h656E;
 buffer[644] = 16'h6167;
 buffer[645] = 16'h6574;
 buffer[646] = 16'h6600;
 buffer[647] = 16'h6147;
 buffer[648] = 16'h6600;
 buffer[649] = 16'h8001;
 buffer[650] = 16'h41AB;
 buffer[651] = 16'h6B8D;
 buffer[652] = 16'h720F;
 buffer[653] = 16'h0504;
 buffer[654] = 16'h2D01;
 buffer[655] = 16'h6D10;
 buffer[656] = 16'h720F;
 buffer[657] = 16'h051C;
 buffer[658] = 16'h6103;
 buffer[659] = 16'h7362;
 buffer[660] = 16'h7A1C;
 buffer[661] = 16'h0524;
 buffer[662] = 16'h6D03;
 buffer[663] = 16'h7861;
 buffer[664] = 16'h7B1F;
 buffer[665] = 16'h052C;
 buffer[666] = 16'h6D03;
 buffer[667] = 16'h6E69;
 buffer[668] = 16'h7C1F;
 buffer[669] = 16'h0534;
 buffer[670] = 16'h7706;
 buffer[671] = 16'h7469;
 buffer[672] = 16'h6968;
 buffer[673] = 16'h006E;
 buffer[674] = 16'h6181;
 buffer[675] = 16'h428F;
 buffer[676] = 16'h6147;
 buffer[677] = 16'h428F;
 buffer[678] = 16'h6B8D;
 buffer[679] = 16'h7F0F;
 buffer[680] = 16'h053C;
 buffer[681] = 16'h7506;
 buffer[682] = 16'h2F6D;
 buffer[683] = 16'h6F6D;
 buffer[684] = 16'h0064;
 buffer[685] = 16'h4279;
 buffer[686] = 16'h6F03;
 buffer[687] = 16'h22D6;
 buffer[688] = 16'h6D10;
 buffer[689] = 16'h800F;
 buffer[690] = 16'h6147;
 buffer[691] = 16'h6147;
 buffer[692] = 16'h6081;
 buffer[693] = 16'h41AB;
 buffer[694] = 16'h6147;
 buffer[695] = 16'h6147;
 buffer[696] = 16'h6081;
 buffer[697] = 16'h41AB;
 buffer[698] = 16'h6B8D;
 buffer[699] = 16'h6203;
 buffer[700] = 16'h6081;
 buffer[701] = 16'h6B8D;
 buffer[702] = 16'h6B81;
 buffer[703] = 16'h6180;
 buffer[704] = 16'h6147;
 buffer[705] = 16'h41AB;
 buffer[706] = 16'h6B8D;
 buffer[707] = 16'h6403;
 buffer[708] = 16'h22CA;
 buffer[709] = 16'h6147;
 buffer[710] = 16'h6103;
 buffer[711] = 16'h6310;
 buffer[712] = 16'h6B8D;
 buffer[713] = 16'h02CB;
 buffer[714] = 16'h6103;
 buffer[715] = 16'h6B8D;
 buffer[716] = 16'h6B81;
 buffer[717] = 16'h22D2;
 buffer[718] = 16'h6B8D;
 buffer[719] = 16'h6A00;
 buffer[720] = 16'h6147;
 buffer[721] = 16'h02B3;
 buffer[722] = 16'h6B8D;
 buffer[723] = 16'h6103;
 buffer[724] = 16'h6103;
 buffer[725] = 16'h718C;
 buffer[726] = 16'h6103;
 buffer[727] = 16'h4273;
 buffer[728] = 16'h8000;
 buffer[729] = 16'h6600;
 buffer[730] = 16'h708D;
 buffer[731] = 16'h0552;
 buffer[732] = 16'h6D05;
 buffer[733] = 16'h6D2F;
 buffer[734] = 16'h646F;
 buffer[735] = 16'h6081;
 buffer[736] = 16'h6810;
 buffer[737] = 16'h6081;
 buffer[738] = 16'h6147;
 buffer[739] = 16'h22E8;
 buffer[740] = 16'h6D10;
 buffer[741] = 16'h6147;
 buffer[742] = 16'h4286;
 buffer[743] = 16'h6B8D;
 buffer[744] = 16'h6147;
 buffer[745] = 16'h6081;
 buffer[746] = 16'h6810;
 buffer[747] = 16'h22EE;
 buffer[748] = 16'h6B81;
 buffer[749] = 16'h6203;
 buffer[750] = 16'h6B8D;
 buffer[751] = 16'h42AD;
 buffer[752] = 16'h6B8D;
 buffer[753] = 16'h22F5;
 buffer[754] = 16'h6180;
 buffer[755] = 16'h6D10;
 buffer[756] = 16'h718C;
 buffer[757] = 16'h700C;
 buffer[758] = 16'h05B8;
 buffer[759] = 16'h2F04;
 buffer[760] = 16'h6F6D;
 buffer[761] = 16'h0064;
 buffer[762] = 16'h6181;
 buffer[763] = 16'h6810;
 buffer[764] = 16'h6180;
 buffer[765] = 16'h02DF;
 buffer[766] = 16'h05EE;
 buffer[767] = 16'h6D03;
 buffer[768] = 16'h646F;
 buffer[769] = 16'h42FA;
 buffer[770] = 16'h710F;
 buffer[771] = 16'h05FE;
 buffer[772] = 16'h2F01;
 buffer[773] = 16'h42FA;
 buffer[774] = 16'h700F;
 buffer[775] = 16'h0608;
 buffer[776] = 16'h7503;
 buffer[777] = 16'h2A6D;
 buffer[778] = 16'h8000;
 buffer[779] = 16'h6180;
 buffer[780] = 16'h800F;
 buffer[781] = 16'h6147;
 buffer[782] = 16'h6081;
 buffer[783] = 16'h41AB;
 buffer[784] = 16'h6147;
 buffer[785] = 16'h6147;
 buffer[786] = 16'h6081;
 buffer[787] = 16'h41AB;
 buffer[788] = 16'h6B8D;
 buffer[789] = 16'h6203;
 buffer[790] = 16'h6B8D;
 buffer[791] = 16'h231D;
 buffer[792] = 16'h6147;
 buffer[793] = 16'h6181;
 buffer[794] = 16'h41AB;
 buffer[795] = 16'h6B8D;
 buffer[796] = 16'h6203;
 buffer[797] = 16'h6B81;
 buffer[798] = 16'h2323;
 buffer[799] = 16'h6B8D;
 buffer[800] = 16'h6A00;
 buffer[801] = 16'h6147;
 buffer[802] = 16'h030E;
 buffer[803] = 16'h6B8D;
 buffer[804] = 16'h6103;
 buffer[805] = 16'h426B;
 buffer[806] = 16'h710F;
 buffer[807] = 16'h0610;
 buffer[808] = 16'h2A01;
 buffer[809] = 16'h430A;
 buffer[810] = 16'h710F;
 buffer[811] = 16'h0650;
 buffer[812] = 16'h6D02;
 buffer[813] = 16'h002A;
 buffer[814] = 16'h4279;
 buffer[815] = 16'h6503;
 buffer[816] = 16'h6810;
 buffer[817] = 16'h6147;
 buffer[818] = 16'h6A10;
 buffer[819] = 16'h6180;
 buffer[820] = 16'h6A10;
 buffer[821] = 16'h430A;
 buffer[822] = 16'h6B8D;
 buffer[823] = 16'h2339;
 buffer[824] = 16'h0286;
 buffer[825] = 16'h700C;
 buffer[826] = 16'h0658;
 buffer[827] = 16'h2A05;
 buffer[828] = 16'h6D2F;
 buffer[829] = 16'h646F;
 buffer[830] = 16'h6147;
 buffer[831] = 16'h432E;
 buffer[832] = 16'h6B8D;
 buffer[833] = 16'h02DF;
 buffer[834] = 16'h0676;
 buffer[835] = 16'h2A02;
 buffer[836] = 16'h002F;
 buffer[837] = 16'h433E;
 buffer[838] = 16'h700F;
 buffer[839] = 16'h0686;
 buffer[840] = 16'h6305;
 buffer[841] = 16'h6C65;
 buffer[842] = 16'h2B6C;
 buffer[843] = 16'h8002;
 buffer[844] = 16'h720F;
 buffer[845] = 16'h0690;
 buffer[846] = 16'h6305;
 buffer[847] = 16'h6C65;
 buffer[848] = 16'h2D6C;
 buffer[849] = 16'h8002;
 buffer[850] = 16'h028F;
 buffer[851] = 16'h069C;
 buffer[852] = 16'h6305;
 buffer[853] = 16'h6C65;
 buffer[854] = 16'h736C;
 buffer[855] = 16'h8001;
 buffer[856] = 16'h7D0F;
 buffer[857] = 16'h06A8;
 buffer[858] = 16'h6202;
 buffer[859] = 16'h006C;
 buffer[860] = 16'h8020;
 buffer[861] = 16'h700C;
 buffer[862] = 16'h06B4;
 buffer[863] = 16'h3E05;
 buffer[864] = 16'h6863;
 buffer[865] = 16'h7261;
 buffer[866] = 16'h807F;
 buffer[867] = 16'h6303;
 buffer[868] = 16'h6081;
 buffer[869] = 16'h807F;
 buffer[870] = 16'h435C;
 buffer[871] = 16'h42A2;
 buffer[872] = 16'h236B;
 buffer[873] = 16'h6103;
 buffer[874] = 16'h805F;
 buffer[875] = 16'h700C;
 buffer[876] = 16'h700C;
 buffer[877] = 16'h06BE;
 buffer[878] = 16'h2B02;
 buffer[879] = 16'h0021;
 buffer[880] = 16'h414F;
 buffer[881] = 16'h6C00;
 buffer[882] = 16'h6203;
 buffer[883] = 16'h6180;
 buffer[884] = 16'h6023;
 buffer[885] = 16'h710F;
 buffer[886] = 16'h06DC;
 buffer[887] = 16'h3202;
 buffer[888] = 16'h0021;
 buffer[889] = 16'h6180;
 buffer[890] = 16'h6181;
 buffer[891] = 16'h6023;
 buffer[892] = 16'h6103;
 buffer[893] = 16'h434B;
 buffer[894] = 16'h6023;
 buffer[895] = 16'h710F;
 buffer[896] = 16'h06EE;
 buffer[897] = 16'h3202;
 buffer[898] = 16'h0040;
 buffer[899] = 16'h6081;
 buffer[900] = 16'h434B;
 buffer[901] = 16'h6C00;
 buffer[902] = 16'h6180;
 buffer[903] = 16'h7C0C;
 buffer[904] = 16'h0702;
 buffer[905] = 16'h6305;
 buffer[906] = 16'h756F;
 buffer[907] = 16'h746E;
 buffer[908] = 16'h6081;
 buffer[909] = 16'h6310;
 buffer[910] = 16'h6180;
 buffer[911] = 16'h017E;
 buffer[912] = 16'h0712;
 buffer[913] = 16'h6804;
 buffer[914] = 16'h7265;
 buffer[915] = 16'h0065;
 buffer[916] = 16'hFEAC;
 buffer[917] = 16'h7C0C;
 buffer[918] = 16'h0722;
 buffer[919] = 16'h6107;
 buffer[920] = 16'h696C;
 buffer[921] = 16'h6E67;
 buffer[922] = 16'h6465;
 buffer[923] = 16'h6081;
 buffer[924] = 16'h8000;
 buffer[925] = 16'h8002;
 buffer[926] = 16'h42AD;
 buffer[927] = 16'h6103;
 buffer[928] = 16'h6081;
 buffer[929] = 16'h23A5;
 buffer[930] = 16'h8002;
 buffer[931] = 16'h6180;
 buffer[932] = 16'h428F;
 buffer[933] = 16'h720F;
 buffer[934] = 16'h072E;
 buffer[935] = 16'h6105;
 buffer[936] = 16'h696C;
 buffer[937] = 16'h6E67;
 buffer[938] = 16'h4394;
 buffer[939] = 16'h439B;
 buffer[940] = 16'hFEAC;
 buffer[941] = 16'h6023;
 buffer[942] = 16'h710F;
 buffer[943] = 16'h074E;
 buffer[944] = 16'h7003;
 buffer[945] = 16'h6461;
 buffer[946] = 16'h4394;
 buffer[947] = 16'h8050;
 buffer[948] = 16'h6203;
 buffer[949] = 16'h039B;
 buffer[950] = 16'h0760;
 buffer[951] = 16'h4008;
 buffer[952] = 16'h7865;
 buffer[953] = 16'h6365;
 buffer[954] = 16'h7475;
 buffer[955] = 16'h0065;
 buffer[956] = 16'h6C00;
 buffer[957] = 16'h4264;
 buffer[958] = 16'h23C0;
 buffer[959] = 16'h0172;
 buffer[960] = 16'h700C;
 buffer[961] = 16'h076E;
 buffer[962] = 16'h6604;
 buffer[963] = 16'h6C69;
 buffer[964] = 16'h006C;
 buffer[965] = 16'h6180;
 buffer[966] = 16'h6147;
 buffer[967] = 16'h6180;
 buffer[968] = 16'h03CC;
 buffer[969] = 16'h4279;
 buffer[970] = 16'h418D;
 buffer[971] = 16'h6310;
 buffer[972] = 16'h6B81;
 buffer[973] = 16'h23D2;
 buffer[974] = 16'h6B8D;
 buffer[975] = 16'h6A00;
 buffer[976] = 16'h6147;
 buffer[977] = 16'h03C9;
 buffer[978] = 16'h6B8D;
 buffer[979] = 16'h6103;
 buffer[980] = 16'h0273;
 buffer[981] = 16'h0784;
 buffer[982] = 16'h6505;
 buffer[983] = 16'h6172;
 buffer[984] = 16'h6573;
 buffer[985] = 16'h8000;
 buffer[986] = 16'h03C5;
 buffer[987] = 16'h07AC;
 buffer[988] = 16'h6405;
 buffer[989] = 16'h6769;
 buffer[990] = 16'h7469;
 buffer[991] = 16'h8009;
 buffer[992] = 16'h6181;
 buffer[993] = 16'h6803;
 buffer[994] = 16'h8007;
 buffer[995] = 16'h6303;
 buffer[996] = 16'h6203;
 buffer[997] = 16'h8030;
 buffer[998] = 16'h720F;
 buffer[999] = 16'h07B8;
 buffer[1000] = 16'h6507;
 buffer[1001] = 16'h7478;
 buffer[1002] = 16'h6172;
 buffer[1003] = 16'h7463;
 buffer[1004] = 16'h8000;
 buffer[1005] = 16'h6180;
 buffer[1006] = 16'h42AD;
 buffer[1007] = 16'h6180;
 buffer[1008] = 16'h03DF;
 buffer[1009] = 16'h07D0;
 buffer[1010] = 16'h3C02;
 buffer[1011] = 16'h0023;
 buffer[1012] = 16'h43B2;
 buffer[1013] = 16'hFE8E;
 buffer[1014] = 16'h6023;
 buffer[1015] = 16'h710F;
 buffer[1016] = 16'h07E4;
 buffer[1017] = 16'h6804;
 buffer[1018] = 16'h6C6F;
 buffer[1019] = 16'h0064;
 buffer[1020] = 16'hFE8E;
 buffer[1021] = 16'h6C00;
 buffer[1022] = 16'h6A00;
 buffer[1023] = 16'h6081;
 buffer[1024] = 16'hFE8E;
 buffer[1025] = 16'h6023;
 buffer[1026] = 16'h6103;
 buffer[1027] = 16'h018D;
 buffer[1028] = 16'h07F2;
 buffer[1029] = 16'h2301;
 buffer[1030] = 16'hFE80;
 buffer[1031] = 16'h6C00;
 buffer[1032] = 16'h43EC;
 buffer[1033] = 16'h03FC;
 buffer[1034] = 16'h080A;
 buffer[1035] = 16'h2302;
 buffer[1036] = 16'h0073;
 buffer[1037] = 16'h4406;
 buffer[1038] = 16'h6081;
 buffer[1039] = 16'h2411;
 buffer[1040] = 16'h040D;
 buffer[1041] = 16'h700C;
 buffer[1042] = 16'h0816;
 buffer[1043] = 16'h7304;
 buffer[1044] = 16'h6769;
 buffer[1045] = 16'h006E;
 buffer[1046] = 16'h6810;
 buffer[1047] = 16'h241A;
 buffer[1048] = 16'h802D;
 buffer[1049] = 16'h03FC;
 buffer[1050] = 16'h700C;
 buffer[1051] = 16'h0826;
 buffer[1052] = 16'h2302;
 buffer[1053] = 16'h003E;
 buffer[1054] = 16'h6103;
 buffer[1055] = 16'hFE8E;
 buffer[1056] = 16'h6C00;
 buffer[1057] = 16'h43B2;
 buffer[1058] = 16'h6181;
 buffer[1059] = 16'h028F;
 buffer[1060] = 16'h0838;
 buffer[1061] = 16'h7303;
 buffer[1062] = 16'h7274;
 buffer[1063] = 16'h6081;
 buffer[1064] = 16'h6147;
 buffer[1065] = 16'h6A10;
 buffer[1066] = 16'h43F4;
 buffer[1067] = 16'h440D;
 buffer[1068] = 16'h6B8D;
 buffer[1069] = 16'h4416;
 buffer[1070] = 16'h041E;
 buffer[1071] = 16'h084A;
 buffer[1072] = 16'h6803;
 buffer[1073] = 16'h7865;
 buffer[1074] = 16'h8010;
 buffer[1075] = 16'hFE80;
 buffer[1076] = 16'h6023;
 buffer[1077] = 16'h710F;
 buffer[1078] = 16'h0860;
 buffer[1079] = 16'h6407;
 buffer[1080] = 16'h6365;
 buffer[1081] = 16'h6D69;
 buffer[1082] = 16'h6C61;
 buffer[1083] = 16'h800A;
 buffer[1084] = 16'hFE80;
 buffer[1085] = 16'h6023;
 buffer[1086] = 16'h710F;
 buffer[1087] = 16'h086E;
 buffer[1088] = 16'h6406;
 buffer[1089] = 16'h6769;
 buffer[1090] = 16'h7469;
 buffer[1091] = 16'h003F;
 buffer[1092] = 16'h6147;
 buffer[1093] = 16'h8030;
 buffer[1094] = 16'h428F;
 buffer[1095] = 16'h8009;
 buffer[1096] = 16'h6181;
 buffer[1097] = 16'h6803;
 buffer[1098] = 16'h2457;
 buffer[1099] = 16'h6081;
 buffer[1100] = 16'h8020;
 buffer[1101] = 16'h6613;
 buffer[1102] = 16'h2451;
 buffer[1103] = 16'h8020;
 buffer[1104] = 16'h428F;
 buffer[1105] = 16'h8007;
 buffer[1106] = 16'h428F;
 buffer[1107] = 16'h6081;
 buffer[1108] = 16'h800A;
 buffer[1109] = 16'h6803;
 buffer[1110] = 16'h6403;
 buffer[1111] = 16'h6081;
 buffer[1112] = 16'h6B8D;
 buffer[1113] = 16'h7F0F;
 buffer[1114] = 16'h0880;
 buffer[1115] = 16'h6E07;
 buffer[1116] = 16'h6D75;
 buffer[1117] = 16'h6562;
 buffer[1118] = 16'h3F72;
 buffer[1119] = 16'hFE80;
 buffer[1120] = 16'h6C00;
 buffer[1121] = 16'h6147;
 buffer[1122] = 16'h8000;
 buffer[1123] = 16'h6181;
 buffer[1124] = 16'h438C;
 buffer[1125] = 16'h6181;
 buffer[1126] = 16'h417E;
 buffer[1127] = 16'h8024;
 buffer[1128] = 16'h6703;
 buffer[1129] = 16'h246F;
 buffer[1130] = 16'h4432;
 buffer[1131] = 16'h6180;
 buffer[1132] = 16'h6310;
 buffer[1133] = 16'h6180;
 buffer[1134] = 16'h6A00;
 buffer[1135] = 16'h6181;
 buffer[1136] = 16'h417E;
 buffer[1137] = 16'h802D;
 buffer[1138] = 16'h6703;
 buffer[1139] = 16'h6147;
 buffer[1140] = 16'h6180;
 buffer[1141] = 16'h6B81;
 buffer[1142] = 16'h428F;
 buffer[1143] = 16'h6180;
 buffer[1144] = 16'h6B81;
 buffer[1145] = 16'h6203;
 buffer[1146] = 16'h4264;
 buffer[1147] = 16'h24A0;
 buffer[1148] = 16'h6A00;
 buffer[1149] = 16'h6147;
 buffer[1150] = 16'h6081;
 buffer[1151] = 16'h6147;
 buffer[1152] = 16'h417E;
 buffer[1153] = 16'hFE80;
 buffer[1154] = 16'h6C00;
 buffer[1155] = 16'h4444;
 buffer[1156] = 16'h249A;
 buffer[1157] = 16'h6180;
 buffer[1158] = 16'hFE80;
 buffer[1159] = 16'h6C00;
 buffer[1160] = 16'h4329;
 buffer[1161] = 16'h6203;
 buffer[1162] = 16'h6B8D;
 buffer[1163] = 16'h6310;
 buffer[1164] = 16'h6B81;
 buffer[1165] = 16'h2492;
 buffer[1166] = 16'h6B8D;
 buffer[1167] = 16'h6A00;
 buffer[1168] = 16'h6147;
 buffer[1169] = 16'h047E;
 buffer[1170] = 16'h6B8D;
 buffer[1171] = 16'h6103;
 buffer[1172] = 16'h6B81;
 buffer[1173] = 16'h6003;
 buffer[1174] = 16'h2498;
 buffer[1175] = 16'h6D10;
 buffer[1176] = 16'h6180;
 buffer[1177] = 16'h049F;
 buffer[1178] = 16'h6B8D;
 buffer[1179] = 16'h6B8D;
 buffer[1180] = 16'h4273;
 buffer[1181] = 16'h4273;
 buffer[1182] = 16'h8000;
 buffer[1183] = 16'h6081;
 buffer[1184] = 16'h6B8D;
 buffer[1185] = 16'h4273;
 buffer[1186] = 16'h6B8D;
 buffer[1187] = 16'hFE80;
 buffer[1188] = 16'h6023;
 buffer[1189] = 16'h710F;
 buffer[1190] = 16'h08B6;
 buffer[1191] = 16'h3F03;
 buffer[1192] = 16'h7872;
 buffer[1193] = 16'h8FFE;
 buffer[1194] = 16'h6600;
 buffer[1195] = 16'h6C00;
 buffer[1196] = 16'h8001;
 buffer[1197] = 16'h6303;
 buffer[1198] = 16'h711C;
 buffer[1199] = 16'h094E;
 buffer[1200] = 16'h7403;
 buffer[1201] = 16'h2178;
 buffer[1202] = 16'h8FFE;
 buffer[1203] = 16'h6600;
 buffer[1204] = 16'h6C00;
 buffer[1205] = 16'h8002;
 buffer[1206] = 16'h6303;
 buffer[1207] = 16'h6010;
 buffer[1208] = 16'h24B2;
 buffer[1209] = 16'h8FFF;
 buffer[1210] = 16'h6600;
 buffer[1211] = 16'h6023;
 buffer[1212] = 16'h710F;
 buffer[1213] = 16'h0960;
 buffer[1214] = 16'h3F04;
 buffer[1215] = 16'h656B;
 buffer[1216] = 16'h0079;
 buffer[1217] = 16'hFEB0;
 buffer[1218] = 16'h03BC;
 buffer[1219] = 16'h097C;
 buffer[1220] = 16'h6504;
 buffer[1221] = 16'h696D;
 buffer[1222] = 16'h0074;
 buffer[1223] = 16'hFEB2;
 buffer[1224] = 16'h03BC;
 buffer[1225] = 16'h0988;
 buffer[1226] = 16'h6B03;
 buffer[1227] = 16'h7965;
 buffer[1228] = 16'h44C1;
 buffer[1229] = 16'h24CC;
 buffer[1230] = 16'h8FFF;
 buffer[1231] = 16'h6600;
 buffer[1232] = 16'h7C0C;
 buffer[1233] = 16'h0994;
 buffer[1234] = 16'h6E04;
 buffer[1235] = 16'h6675;
 buffer[1236] = 16'h003F;
 buffer[1237] = 16'h44C1;
 buffer[1238] = 16'h6081;
 buffer[1239] = 16'h24DC;
 buffer[1240] = 16'h6103;
 buffer[1241] = 16'h44CC;
 buffer[1242] = 16'h800D;
 buffer[1243] = 16'h770F;
 buffer[1244] = 16'h700C;
 buffer[1245] = 16'h09A4;
 buffer[1246] = 16'h7406;
 buffer[1247] = 16'h6D69;
 buffer[1248] = 16'h7265;
 buffer[1249] = 16'h0040;
 buffer[1250] = 16'h8FFB;
 buffer[1251] = 16'h6600;
 buffer[1252] = 16'h7C0C;
 buffer[1253] = 16'h09BC;
 buffer[1254] = 16'h6C04;
 buffer[1255] = 16'h6465;
 buffer[1256] = 16'h0040;
 buffer[1257] = 16'h8FFD;
 buffer[1258] = 16'h6600;
 buffer[1259] = 16'h7C0C;
 buffer[1260] = 16'h09CC;
 buffer[1261] = 16'h6C04;
 buffer[1262] = 16'h6465;
 buffer[1263] = 16'h0021;
 buffer[1264] = 16'h8FFD;
 buffer[1265] = 16'h6600;
 buffer[1266] = 16'h6023;
 buffer[1267] = 16'h710F;
 buffer[1268] = 16'h09DA;
 buffer[1269] = 16'h6208;
 buffer[1270] = 16'h7475;
 buffer[1271] = 16'h6F74;
 buffer[1272] = 16'h736E;
 buffer[1273] = 16'h0040;
 buffer[1274] = 16'h8FFC;
 buffer[1275] = 16'h6600;
 buffer[1276] = 16'h7C0C;
 buffer[1277] = 16'h09EA;
 buffer[1278] = 16'h7305;
 buffer[1279] = 16'h6170;
 buffer[1280] = 16'h6563;
 buffer[1281] = 16'h435C;
 buffer[1282] = 16'h04C7;
 buffer[1283] = 16'h09FC;
 buffer[1284] = 16'h7306;
 buffer[1285] = 16'h6170;
 buffer[1286] = 16'h6563;
 buffer[1287] = 16'h0073;
 buffer[1288] = 16'h8000;
 buffer[1289] = 16'h6B13;
 buffer[1290] = 16'h6147;
 buffer[1291] = 16'h050D;
 buffer[1292] = 16'h4501;
 buffer[1293] = 16'h6B81;
 buffer[1294] = 16'h2513;
 buffer[1295] = 16'h6B8D;
 buffer[1296] = 16'h6A00;
 buffer[1297] = 16'h6147;
 buffer[1298] = 16'h050C;
 buffer[1299] = 16'h6B8D;
 buffer[1300] = 16'h710F;
 buffer[1301] = 16'h0A08;
 buffer[1302] = 16'h7404;
 buffer[1303] = 16'h7079;
 buffer[1304] = 16'h0065;
 buffer[1305] = 16'h6147;
 buffer[1306] = 16'h051D;
 buffer[1307] = 16'h438C;
 buffer[1308] = 16'h44C7;
 buffer[1309] = 16'h6B81;
 buffer[1310] = 16'h2523;
 buffer[1311] = 16'h6B8D;
 buffer[1312] = 16'h6A00;
 buffer[1313] = 16'h6147;
 buffer[1314] = 16'h051B;
 buffer[1315] = 16'h6B8D;
 buffer[1316] = 16'h6103;
 buffer[1317] = 16'h710F;
 buffer[1318] = 16'h0A2C;
 buffer[1319] = 16'h6302;
 buffer[1320] = 16'h0072;
 buffer[1321] = 16'h800D;
 buffer[1322] = 16'h44C7;
 buffer[1323] = 16'h800A;
 buffer[1324] = 16'h04C7;
 buffer[1325] = 16'h0A4E;
 buffer[1326] = 16'h6443;
 buffer[1327] = 16'h246F;
 buffer[1328] = 16'h6B8D;
 buffer[1329] = 16'h6B81;
 buffer[1330] = 16'h6B8D;
 buffer[1331] = 16'h438C;
 buffer[1332] = 16'h6203;
 buffer[1333] = 16'h439B;
 buffer[1334] = 16'h6147;
 buffer[1335] = 16'h6180;
 buffer[1336] = 16'h6147;
 buffer[1337] = 16'h700C;
 buffer[1338] = 16'h0A5C;
 buffer[1339] = 16'h2443;
 buffer[1340] = 16'h7C22;
 buffer[1341] = 16'h4530;
 buffer[1342] = 16'h700C;
 buffer[1343] = 16'h0A76;
 buffer[1344] = 16'h2E02;
 buffer[1345] = 16'h0024;
 buffer[1346] = 16'h438C;
 buffer[1347] = 16'h0519;
 buffer[1348] = 16'h0A80;
 buffer[1349] = 16'h2E43;
 buffer[1350] = 16'h7C22;
 buffer[1351] = 16'h4530;
 buffer[1352] = 16'h0542;
 buffer[1353] = 16'h0A8A;
 buffer[1354] = 16'h2E02;
 buffer[1355] = 16'h0072;
 buffer[1356] = 16'h6147;
 buffer[1357] = 16'h4427;
 buffer[1358] = 16'h6B8D;
 buffer[1359] = 16'h6181;
 buffer[1360] = 16'h428F;
 buffer[1361] = 16'h4508;
 buffer[1362] = 16'h0519;
 buffer[1363] = 16'h0A94;
 buffer[1364] = 16'h7503;
 buffer[1365] = 16'h722E;
 buffer[1366] = 16'h6147;
 buffer[1367] = 16'h43F4;
 buffer[1368] = 16'h440D;
 buffer[1369] = 16'h441E;
 buffer[1370] = 16'h6B8D;
 buffer[1371] = 16'h6181;
 buffer[1372] = 16'h428F;
 buffer[1373] = 16'h4508;
 buffer[1374] = 16'h0519;
 buffer[1375] = 16'h0AA8;
 buffer[1376] = 16'h7502;
 buffer[1377] = 16'h002E;
 buffer[1378] = 16'h43F4;
 buffer[1379] = 16'h440D;
 buffer[1380] = 16'h441E;
 buffer[1381] = 16'h4501;
 buffer[1382] = 16'h0519;
 buffer[1383] = 16'h0AC0;
 buffer[1384] = 16'h2E01;
 buffer[1385] = 16'hFE80;
 buffer[1386] = 16'h6C00;
 buffer[1387] = 16'h800A;
 buffer[1388] = 16'h6503;
 buffer[1389] = 16'h256F;
 buffer[1390] = 16'h0562;
 buffer[1391] = 16'h4427;
 buffer[1392] = 16'h4501;
 buffer[1393] = 16'h0519;
 buffer[1394] = 16'h0AD0;
 buffer[1395] = 16'h2E02;
 buffer[1396] = 16'h0023;
 buffer[1397] = 16'hFE80;
 buffer[1398] = 16'h6C00;
 buffer[1399] = 16'h6180;
 buffer[1400] = 16'h443B;
 buffer[1401] = 16'h4569;
 buffer[1402] = 16'hFE80;
 buffer[1403] = 16'h6023;
 buffer[1404] = 16'h710F;
 buffer[1405] = 16'h0AE6;
 buffer[1406] = 16'h7503;
 buffer[1407] = 16'h232E;
 buffer[1408] = 16'hFE80;
 buffer[1409] = 16'h6C00;
 buffer[1410] = 16'h6180;
 buffer[1411] = 16'h443B;
 buffer[1412] = 16'h43F4;
 buffer[1413] = 16'h440D;
 buffer[1414] = 16'h441E;
 buffer[1415] = 16'h4501;
 buffer[1416] = 16'h4519;
 buffer[1417] = 16'hFE80;
 buffer[1418] = 16'h6023;
 buffer[1419] = 16'h710F;
 buffer[1420] = 16'h0AFC;
 buffer[1421] = 16'h7504;
 buffer[1422] = 16'h722E;
 buffer[1423] = 16'h0023;
 buffer[1424] = 16'hFE80;
 buffer[1425] = 16'h6C00;
 buffer[1426] = 16'h426B;
 buffer[1427] = 16'h426B;
 buffer[1428] = 16'h443B;
 buffer[1429] = 16'h6147;
 buffer[1430] = 16'h43F4;
 buffer[1431] = 16'h440D;
 buffer[1432] = 16'h441E;
 buffer[1433] = 16'h6B8D;
 buffer[1434] = 16'h6181;
 buffer[1435] = 16'h428F;
 buffer[1436] = 16'h4508;
 buffer[1437] = 16'h4519;
 buffer[1438] = 16'hFE80;
 buffer[1439] = 16'h6023;
 buffer[1440] = 16'h710F;
 buffer[1441] = 16'h0B1A;
 buffer[1442] = 16'h2E03;
 buffer[1443] = 16'h2372;
 buffer[1444] = 16'hFE80;
 buffer[1445] = 16'h6C00;
 buffer[1446] = 16'h426B;
 buffer[1447] = 16'h426B;
 buffer[1448] = 16'h443B;
 buffer[1449] = 16'h6147;
 buffer[1450] = 16'h4427;
 buffer[1451] = 16'h6B8D;
 buffer[1452] = 16'h6181;
 buffer[1453] = 16'h428F;
 buffer[1454] = 16'h4508;
 buffer[1455] = 16'h4519;
 buffer[1456] = 16'hFE80;
 buffer[1457] = 16'h6023;
 buffer[1458] = 16'h710F;
 buffer[1459] = 16'h0B44;
 buffer[1460] = 16'h6305;
 buffer[1461] = 16'h6F6D;
 buffer[1462] = 16'h6576;
 buffer[1463] = 16'h6147;
 buffer[1464] = 16'h05C1;
 buffer[1465] = 16'h6147;
 buffer[1466] = 16'h6081;
 buffer[1467] = 16'h417E;
 buffer[1468] = 16'h6B81;
 buffer[1469] = 16'h418D;
 buffer[1470] = 16'h6310;
 buffer[1471] = 16'h6B8D;
 buffer[1472] = 16'h6310;
 buffer[1473] = 16'h6B81;
 buffer[1474] = 16'h25C7;
 buffer[1475] = 16'h6B8D;
 buffer[1476] = 16'h6A00;
 buffer[1477] = 16'h6147;
 buffer[1478] = 16'h05B9;
 buffer[1479] = 16'h6B8D;
 buffer[1480] = 16'h6103;
 buffer[1481] = 16'h0273;
 buffer[1482] = 16'h0B68;
 buffer[1483] = 16'h7005;
 buffer[1484] = 16'h6361;
 buffer[1485] = 16'h246B;
 buffer[1486] = 16'h6081;
 buffer[1487] = 16'h6147;
 buffer[1488] = 16'h4279;
 buffer[1489] = 16'h6023;
 buffer[1490] = 16'h6103;
 buffer[1491] = 16'h6310;
 buffer[1492] = 16'h6180;
 buffer[1493] = 16'h45B7;
 buffer[1494] = 16'h6B8D;
 buffer[1495] = 16'h700C;
 buffer[1496] = 16'h0B96;
 buffer[1497] = 16'h3F01;
 buffer[1498] = 16'h6C00;
 buffer[1499] = 16'h0569;
 buffer[1500] = 16'h0BB2;
 buffer[1501] = 16'h3205;
 buffer[1502] = 16'h766F;
 buffer[1503] = 16'h7265;
 buffer[1504] = 16'h6147;
 buffer[1505] = 16'h6147;
 buffer[1506] = 16'h4279;
 buffer[1507] = 16'h6B8D;
 buffer[1508] = 16'h6B8D;
 buffer[1509] = 16'h426B;
 buffer[1510] = 16'h6147;
 buffer[1511] = 16'h426B;
 buffer[1512] = 16'h6B8D;
 buffer[1513] = 16'h700C;
 buffer[1514] = 16'h0BBA;
 buffer[1515] = 16'h3205;
 buffer[1516] = 16'h7773;
 buffer[1517] = 16'h7061;
 buffer[1518] = 16'h426B;
 buffer[1519] = 16'h6147;
 buffer[1520] = 16'h426B;
 buffer[1521] = 16'h6B8D;
 buffer[1522] = 16'h700C;
 buffer[1523] = 16'h0BD6;
 buffer[1524] = 16'h3204;
 buffer[1525] = 16'h696E;
 buffer[1526] = 16'h0070;
 buffer[1527] = 16'h426B;
 buffer[1528] = 16'h6103;
 buffer[1529] = 16'h426B;
 buffer[1530] = 16'h710F;
 buffer[1531] = 16'h0BE8;
 buffer[1532] = 16'h3204;
 buffer[1533] = 16'h6F72;
 buffer[1534] = 16'h0074;
 buffer[1535] = 16'h6180;
 buffer[1536] = 16'h6147;
 buffer[1537] = 16'h6147;
 buffer[1538] = 16'h45EE;
 buffer[1539] = 16'h6B8D;
 buffer[1540] = 16'h6B8D;
 buffer[1541] = 16'h6180;
 buffer[1542] = 16'h05EE;
 buffer[1543] = 16'h0BF8;
 buffer[1544] = 16'h6402;
 buffer[1545] = 16'h003D;
 buffer[1546] = 16'h6147;
 buffer[1547] = 16'h426B;
 buffer[1548] = 16'h6503;
 buffer[1549] = 16'h6180;
 buffer[1550] = 16'h6B8D;
 buffer[1551] = 16'h6503;
 buffer[1552] = 16'h6403;
 buffer[1553] = 16'h701C;
 buffer[1554] = 16'h0C10;
 buffer[1555] = 16'h6403;
 buffer[1556] = 16'h3E3C;
 buffer[1557] = 16'h460A;
 buffer[1558] = 16'h760C;
 buffer[1559] = 16'h0C26;
 buffer[1560] = 16'h6402;
 buffer[1561] = 16'h002B;
 buffer[1562] = 16'h426B;
 buffer[1563] = 16'h6203;
 buffer[1564] = 16'h6147;
 buffer[1565] = 16'h6181;
 buffer[1566] = 16'h6203;
 buffer[1567] = 16'h6081;
 buffer[1568] = 16'h426B;
 buffer[1569] = 16'h6F03;
 buffer[1570] = 16'h2626;
 buffer[1571] = 16'h6B8D;
 buffer[1572] = 16'h6310;
 buffer[1573] = 16'h0627;
 buffer[1574] = 16'h6B8D;
 buffer[1575] = 16'h700C;
 buffer[1576] = 16'h0C30;
 buffer[1577] = 16'h6402;
 buffer[1578] = 16'h002D;
 buffer[1579] = 16'h4286;
 buffer[1580] = 16'h061A;
 buffer[1581] = 16'h0C52;
 buffer[1582] = 16'h7303;
 buffer[1583] = 16'h643E;
 buffer[1584] = 16'h6081;
 buffer[1585] = 16'h781C;
 buffer[1586] = 16'h0C5C;
 buffer[1587] = 16'h6403;
 buffer[1588] = 16'h2B31;
 buffer[1589] = 16'h8001;
 buffer[1590] = 16'h4630;
 buffer[1591] = 16'h061A;
 buffer[1592] = 16'h0C66;
 buffer[1593] = 16'h6404;
 buffer[1594] = 16'h6F78;
 buffer[1595] = 16'h0072;
 buffer[1596] = 16'h426B;
 buffer[1597] = 16'h6503;
 buffer[1598] = 16'h4155;
 buffer[1599] = 16'h6503;
 buffer[1600] = 16'h718C;
 buffer[1601] = 16'h0C72;
 buffer[1602] = 16'h6404;
 buffer[1603] = 16'h6E61;
 buffer[1604] = 16'h0064;
 buffer[1605] = 16'h426B;
 buffer[1606] = 16'h6303;
 buffer[1607] = 16'h4155;
 buffer[1608] = 16'h6303;
 buffer[1609] = 16'h718C;
 buffer[1610] = 16'h0C84;
 buffer[1611] = 16'h6403;
 buffer[1612] = 16'h726F;
 buffer[1613] = 16'h426B;
 buffer[1614] = 16'h6403;
 buffer[1615] = 16'h4155;
 buffer[1616] = 16'h6403;
 buffer[1617] = 16'h718C;
 buffer[1618] = 16'h0C96;
 buffer[1619] = 16'h6407;
 buffer[1620] = 16'h6E69;
 buffer[1621] = 16'h6576;
 buffer[1622] = 16'h7472;
 buffer[1623] = 16'h6600;
 buffer[1624] = 16'h6180;
 buffer[1625] = 16'h6600;
 buffer[1626] = 16'h718C;
 buffer[1627] = 16'h0CA6;
 buffer[1628] = 16'h6402;
 buffer[1629] = 16'h003C;
 buffer[1630] = 16'h426B;
 buffer[1631] = 16'h4279;
 buffer[1632] = 16'h6703;
 buffer[1633] = 16'h2665;
 buffer[1634] = 16'h4273;
 buffer[1635] = 16'h6F03;
 buffer[1636] = 16'h0667;
 buffer[1637] = 16'h45F7;
 buffer[1638] = 16'h761F;
 buffer[1639] = 16'h0CB8;
 buffer[1640] = 16'h6402;
 buffer[1641] = 16'h003E;
 buffer[1642] = 16'h45EE;
 buffer[1643] = 16'h065E;
 buffer[1644] = 16'h0CD0;
 buffer[1645] = 16'h6403;
 buffer[1646] = 16'h3D30;
 buffer[1647] = 16'h6403;
 buffer[1648] = 16'h701C;
 buffer[1649] = 16'h0CDA;
 buffer[1650] = 16'h6403;
 buffer[1651] = 16'h3C30;
 buffer[1652] = 16'h8000;
 buffer[1653] = 16'h4630;
 buffer[1654] = 16'h065E;
 buffer[1655] = 16'h0CE4;
 buffer[1656] = 16'h6404;
 buffer[1657] = 16'h3C30;
 buffer[1658] = 16'h003E;
 buffer[1659] = 16'h466F;
 buffer[1660] = 16'h760C;
 buffer[1661] = 16'h0CF0;
 buffer[1662] = 16'h6403;
 buffer[1663] = 16'h2A32;
 buffer[1664] = 16'h4279;
 buffer[1665] = 16'h061A;
 buffer[1666] = 16'h0CFC;
 buffer[1667] = 16'h6403;
 buffer[1668] = 16'h2F32;
 buffer[1669] = 16'h6081;
 buffer[1670] = 16'h800F;
 buffer[1671] = 16'h6D03;
 buffer[1672] = 16'h6147;
 buffer[1673] = 16'h415D;
 buffer[1674] = 16'h6180;
 buffer[1675] = 16'h415D;
 buffer[1676] = 16'h6B8D;
 buffer[1677] = 16'h6403;
 buffer[1678] = 16'h718C;
 buffer[1679] = 16'h0D06;
 buffer[1680] = 16'h6403;
 buffer[1681] = 16'h2D31;
 buffer[1682] = 16'h8001;
 buffer[1683] = 16'h4630;
 buffer[1684] = 16'h4286;
 buffer[1685] = 16'h061A;
 buffer[1686] = 16'h0D20;
 buffer[1687] = 16'h7308;
 buffer[1688] = 16'h7465;
 buffer[1689] = 16'h6970;
 buffer[1690] = 16'h6578;
 buffer[1691] = 16'h006C;
 buffer[1692] = 16'h80FE;
 buffer[1693] = 16'h6600;
 buffer[1694] = 16'h6023;
 buffer[1695] = 16'h6103;
 buffer[1696] = 16'h80FF;
 buffer[1697] = 16'h6600;
 buffer[1698] = 16'h6023;
 buffer[1699] = 16'h6103;
 buffer[1700] = 16'h80FD;
 buffer[1701] = 16'h6600;
 buffer[1702] = 16'h6023;
 buffer[1703] = 16'h710F;
 buffer[1704] = 16'h0D2E;
 buffer[1705] = 16'h7307;
 buffer[1706] = 16'h7465;
 buffer[1707] = 16'h6863;
 buffer[1708] = 16'h7261;
 buffer[1709] = 16'h80EE;
 buffer[1710] = 16'h6600;
 buffer[1711] = 16'h6023;
 buffer[1712] = 16'h6103;
 buffer[1713] = 16'h80EF;
 buffer[1714] = 16'h6600;
 buffer[1715] = 16'h6023;
 buffer[1716] = 16'h6103;
 buffer[1717] = 16'h80EC;
 buffer[1718] = 16'h6600;
 buffer[1719] = 16'h6023;
 buffer[1720] = 16'h6103;
 buffer[1721] = 16'h80EB;
 buffer[1722] = 16'h6600;
 buffer[1723] = 16'h6023;
 buffer[1724] = 16'h6103;
 buffer[1725] = 16'h80ED;
 buffer[1726] = 16'h6600;
 buffer[1727] = 16'h6023;
 buffer[1728] = 16'h710F;
 buffer[1729] = 16'h0D52;
 buffer[1730] = 16'h2807;
 buffer[1731] = 16'h6170;
 buffer[1732] = 16'h7372;
 buffer[1733] = 16'h2965;
 buffer[1734] = 16'hFE82;
 buffer[1735] = 16'h6023;
 buffer[1736] = 16'h6103;
 buffer[1737] = 16'h6181;
 buffer[1738] = 16'h6147;
 buffer[1739] = 16'h6081;
 buffer[1740] = 16'h2711;
 buffer[1741] = 16'h6A00;
 buffer[1742] = 16'hFE82;
 buffer[1743] = 16'h6C00;
 buffer[1744] = 16'h435C;
 buffer[1745] = 16'h6703;
 buffer[1746] = 16'h26ED;
 buffer[1747] = 16'h6147;
 buffer[1748] = 16'h438C;
 buffer[1749] = 16'hFE82;
 buffer[1750] = 16'h6C00;
 buffer[1751] = 16'h6180;
 buffer[1752] = 16'h428F;
 buffer[1753] = 16'h6810;
 buffer[1754] = 16'h6600;
 buffer[1755] = 16'h6B81;
 buffer[1756] = 16'h6910;
 buffer[1757] = 16'h6303;
 buffer[1758] = 16'h26EB;
 buffer[1759] = 16'h6B81;
 buffer[1760] = 16'h26E5;
 buffer[1761] = 16'h6B8D;
 buffer[1762] = 16'h6A00;
 buffer[1763] = 16'h6147;
 buffer[1764] = 16'h06D4;
 buffer[1765] = 16'h6B8D;
 buffer[1766] = 16'h6103;
 buffer[1767] = 16'h6B8D;
 buffer[1768] = 16'h6103;
 buffer[1769] = 16'h8000;
 buffer[1770] = 16'h708D;
 buffer[1771] = 16'h6A00;
 buffer[1772] = 16'h6B8D;
 buffer[1773] = 16'h6181;
 buffer[1774] = 16'h6180;
 buffer[1775] = 16'h6147;
 buffer[1776] = 16'h438C;
 buffer[1777] = 16'hFE82;
 buffer[1778] = 16'h6C00;
 buffer[1779] = 16'h6180;
 buffer[1780] = 16'h428F;
 buffer[1781] = 16'hFE82;
 buffer[1782] = 16'h6C00;
 buffer[1783] = 16'h435C;
 buffer[1784] = 16'h6703;
 buffer[1785] = 16'h26FB;
 buffer[1786] = 16'h6810;
 buffer[1787] = 16'h2707;
 buffer[1788] = 16'h6B81;
 buffer[1789] = 16'h2702;
 buffer[1790] = 16'h6B8D;
 buffer[1791] = 16'h6A00;
 buffer[1792] = 16'h6147;
 buffer[1793] = 16'h06F0;
 buffer[1794] = 16'h6B8D;
 buffer[1795] = 16'h6103;
 buffer[1796] = 16'h6081;
 buffer[1797] = 16'h6147;
 buffer[1798] = 16'h070C;
 buffer[1799] = 16'h6B8D;
 buffer[1800] = 16'h6103;
 buffer[1801] = 16'h6081;
 buffer[1802] = 16'h6147;
 buffer[1803] = 16'h6A00;
 buffer[1804] = 16'h6181;
 buffer[1805] = 16'h428F;
 buffer[1806] = 16'h6B8D;
 buffer[1807] = 16'h6B8D;
 buffer[1808] = 16'h028F;
 buffer[1809] = 16'h6181;
 buffer[1810] = 16'h6B8D;
 buffer[1811] = 16'h028F;
 buffer[1812] = 16'h0D84;
 buffer[1813] = 16'h7005;
 buffer[1814] = 16'h7261;
 buffer[1815] = 16'h6573;
 buffer[1816] = 16'h6147;
 buffer[1817] = 16'hFE88;
 buffer[1818] = 16'h6C00;
 buffer[1819] = 16'hFE84;
 buffer[1820] = 16'h6C00;
 buffer[1821] = 16'h6203;
 buffer[1822] = 16'hFE86;
 buffer[1823] = 16'h6C00;
 buffer[1824] = 16'hFE84;
 buffer[1825] = 16'h6C00;
 buffer[1826] = 16'h428F;
 buffer[1827] = 16'h6B8D;
 buffer[1828] = 16'h46C6;
 buffer[1829] = 16'hFE84;
 buffer[1830] = 16'h0370;
 buffer[1831] = 16'h0E2A;
 buffer[1832] = 16'h2E82;
 buffer[1833] = 16'h0028;
 buffer[1834] = 16'h8029;
 buffer[1835] = 16'h4718;
 buffer[1836] = 16'h0519;
 buffer[1837] = 16'h0E50;
 buffer[1838] = 16'h2881;
 buffer[1839] = 16'h8029;
 buffer[1840] = 16'h4718;
 buffer[1841] = 16'h0273;
 buffer[1842] = 16'h0E5C;
 buffer[1843] = 16'h3C83;
 buffer[1844] = 16'h3E5C;
 buffer[1845] = 16'hFE86;
 buffer[1846] = 16'h6C00;
 buffer[1847] = 16'hFE84;
 buffer[1848] = 16'h6023;
 buffer[1849] = 16'h710F;
 buffer[1850] = 16'h0E66;
 buffer[1851] = 16'h5C81;
 buffer[1852] = 16'hFEB6;
 buffer[1853] = 16'h03BC;
 buffer[1854] = 16'h0E76;
 buffer[1855] = 16'h7704;
 buffer[1856] = 16'h726F;
 buffer[1857] = 16'h0064;
 buffer[1858] = 16'h4718;
 buffer[1859] = 16'h4394;
 buffer[1860] = 16'h434B;
 buffer[1861] = 16'h05CE;
 buffer[1862] = 16'h0E7E;
 buffer[1863] = 16'h7405;
 buffer[1864] = 16'h6B6F;
 buffer[1865] = 16'h6E65;
 buffer[1866] = 16'h435C;
 buffer[1867] = 16'h0742;
 buffer[1868] = 16'h0E8E;
 buffer[1869] = 16'h6E05;
 buffer[1870] = 16'h6D61;
 buffer[1871] = 16'h3E65;
 buffer[1872] = 16'h438C;
 buffer[1873] = 16'h801F;
 buffer[1874] = 16'h6303;
 buffer[1875] = 16'h6203;
 buffer[1876] = 16'h039B;
 buffer[1877] = 16'h0E9A;
 buffer[1878] = 16'h7305;
 buffer[1879] = 16'h6D61;
 buffer[1880] = 16'h3F65;
 buffer[1881] = 16'h6A00;
 buffer[1882] = 16'h6147;
 buffer[1883] = 16'h0769;
 buffer[1884] = 16'h6181;
 buffer[1885] = 16'h6B81;
 buffer[1886] = 16'h6203;
 buffer[1887] = 16'h417E;
 buffer[1888] = 16'h6181;
 buffer[1889] = 16'h6B81;
 buffer[1890] = 16'h6203;
 buffer[1891] = 16'h417E;
 buffer[1892] = 16'h428F;
 buffer[1893] = 16'h4264;
 buffer[1894] = 16'h2769;
 buffer[1895] = 16'h6B8D;
 buffer[1896] = 16'h710F;
 buffer[1897] = 16'h6B81;
 buffer[1898] = 16'h276F;
 buffer[1899] = 16'h6B8D;
 buffer[1900] = 16'h6A00;
 buffer[1901] = 16'h6147;
 buffer[1902] = 16'h075C;
 buffer[1903] = 16'h6B8D;
 buffer[1904] = 16'h6103;
 buffer[1905] = 16'h8000;
 buffer[1906] = 16'h700C;
 buffer[1907] = 16'h0EAC;
 buffer[1908] = 16'h6604;
 buffer[1909] = 16'h6E69;
 buffer[1910] = 16'h0064;
 buffer[1911] = 16'h6180;
 buffer[1912] = 16'h6081;
 buffer[1913] = 16'h417E;
 buffer[1914] = 16'hFE82;
 buffer[1915] = 16'h6023;
 buffer[1916] = 16'h6103;
 buffer[1917] = 16'h6081;
 buffer[1918] = 16'h6C00;
 buffer[1919] = 16'h6147;
 buffer[1920] = 16'h434B;
 buffer[1921] = 16'h6180;
 buffer[1922] = 16'h6C00;
 buffer[1923] = 16'h6081;
 buffer[1924] = 16'h2795;
 buffer[1925] = 16'h6081;
 buffer[1926] = 16'h6C00;
 buffer[1927] = 16'hFF1F;
 buffer[1928] = 16'h6303;
 buffer[1929] = 16'h6B81;
 buffer[1930] = 16'h6503;
 buffer[1931] = 16'h2790;
 buffer[1932] = 16'h434B;
 buffer[1933] = 16'h8000;
 buffer[1934] = 16'h6600;
 buffer[1935] = 16'h0794;
 buffer[1936] = 16'h434B;
 buffer[1937] = 16'hFE82;
 buffer[1938] = 16'h6C00;
 buffer[1939] = 16'h4759;
 buffer[1940] = 16'h079A;
 buffer[1941] = 16'h6B8D;
 buffer[1942] = 16'h6103;
 buffer[1943] = 16'h6180;
 buffer[1944] = 16'h4351;
 buffer[1945] = 16'h718C;
 buffer[1946] = 16'h279F;
 buffer[1947] = 16'h8002;
 buffer[1948] = 16'h4357;
 buffer[1949] = 16'h428F;
 buffer[1950] = 16'h0782;
 buffer[1951] = 16'h6B8D;
 buffer[1952] = 16'h6103;
 buffer[1953] = 16'h6003;
 buffer[1954] = 16'h4351;
 buffer[1955] = 16'h6081;
 buffer[1956] = 16'h4750;
 buffer[1957] = 16'h718C;
 buffer[1958] = 16'h0EE8;
 buffer[1959] = 16'h3C07;
 buffer[1960] = 16'h616E;
 buffer[1961] = 16'h656D;
 buffer[1962] = 16'h3E3F;
 buffer[1963] = 16'hFE90;
 buffer[1964] = 16'h6081;
 buffer[1965] = 16'h4383;
 buffer[1966] = 16'h6503;
 buffer[1967] = 16'h27B1;
 buffer[1968] = 16'h4351;
 buffer[1969] = 16'h6147;
 buffer[1970] = 16'h6B8D;
 buffer[1971] = 16'h434B;
 buffer[1972] = 16'h6081;
 buffer[1973] = 16'h6147;
 buffer[1974] = 16'h6C00;
 buffer[1975] = 16'h4264;
 buffer[1976] = 16'h27BE;
 buffer[1977] = 16'h4777;
 buffer[1978] = 16'h4264;
 buffer[1979] = 16'h27B2;
 buffer[1980] = 16'h6B8D;
 buffer[1981] = 16'h710F;
 buffer[1982] = 16'h6B8D;
 buffer[1983] = 16'h6103;
 buffer[1984] = 16'h8000;
 buffer[1985] = 16'h700C;
 buffer[1986] = 16'h0F4E;
 buffer[1987] = 16'h6E05;
 buffer[1988] = 16'h6D61;
 buffer[1989] = 16'h3F65;
 buffer[1990] = 16'hFEB8;
 buffer[1991] = 16'h03BC;
 buffer[1992] = 16'h0F86;
 buffer[1993] = 16'h5E02;
 buffer[1994] = 16'h0068;
 buffer[1995] = 16'h6147;
 buffer[1996] = 16'h6181;
 buffer[1997] = 16'h6B81;
 buffer[1998] = 16'h6803;
 buffer[1999] = 16'h6081;
 buffer[2000] = 16'h27D6;
 buffer[2001] = 16'h8008;
 buffer[2002] = 16'h6081;
 buffer[2003] = 16'h44C7;
 buffer[2004] = 16'h4501;
 buffer[2005] = 16'h44C7;
 buffer[2006] = 16'h6B8D;
 buffer[2007] = 16'h720F;
 buffer[2008] = 16'h0F92;
 buffer[2009] = 16'h7403;
 buffer[2010] = 16'h7061;
 buffer[2011] = 16'h6081;
 buffer[2012] = 16'h44C7;
 buffer[2013] = 16'h6181;
 buffer[2014] = 16'h418D;
 buffer[2015] = 16'h731C;
 buffer[2016] = 16'h0FB2;
 buffer[2017] = 16'h6B04;
 buffer[2018] = 16'h6174;
 buffer[2019] = 16'h0070;
 buffer[2020] = 16'h6081;
 buffer[2021] = 16'h800D;
 buffer[2022] = 16'h6503;
 buffer[2023] = 16'h27EE;
 buffer[2024] = 16'h8008;
 buffer[2025] = 16'h6503;
 buffer[2026] = 16'h27ED;
 buffer[2027] = 16'h435C;
 buffer[2028] = 16'h07DB;
 buffer[2029] = 16'h07CB;
 buffer[2030] = 16'h6103;
 buffer[2031] = 16'h6003;
 buffer[2032] = 16'h708D;
 buffer[2033] = 16'h0FC2;
 buffer[2034] = 16'h6106;
 buffer[2035] = 16'h6363;
 buffer[2036] = 16'h7065;
 buffer[2037] = 16'h0074;
 buffer[2038] = 16'h6181;
 buffer[2039] = 16'h6203;
 buffer[2040] = 16'h6181;
 buffer[2041] = 16'h4279;
 buffer[2042] = 16'h6503;
 buffer[2043] = 16'h2807;
 buffer[2044] = 16'h44CC;
 buffer[2045] = 16'h6081;
 buffer[2046] = 16'h435C;
 buffer[2047] = 16'h428F;
 buffer[2048] = 16'h807F;
 buffer[2049] = 16'h6F03;
 buffer[2050] = 16'h2805;
 buffer[2051] = 16'h47DB;
 buffer[2052] = 16'h0806;
 buffer[2053] = 16'h47E4;
 buffer[2054] = 16'h07F9;
 buffer[2055] = 16'h6103;
 buffer[2056] = 16'h6181;
 buffer[2057] = 16'h028F;
 buffer[2058] = 16'h0FE4;
 buffer[2059] = 16'h7105;
 buffer[2060] = 16'h6575;
 buffer[2061] = 16'h7972;
 buffer[2062] = 16'hFE88;
 buffer[2063] = 16'h6C00;
 buffer[2064] = 16'h8050;
 buffer[2065] = 16'h47F6;
 buffer[2066] = 16'hFE86;
 buffer[2067] = 16'h6023;
 buffer[2068] = 16'h6103;
 buffer[2069] = 16'h6103;
 buffer[2070] = 16'h8000;
 buffer[2071] = 16'hFE84;
 buffer[2072] = 16'h6023;
 buffer[2073] = 16'h710F;
 buffer[2074] = 16'h1016;
 buffer[2075] = 16'h6106;
 buffer[2076] = 16'h6F62;
 buffer[2077] = 16'h7472;
 buffer[2078] = 16'h0032;
 buffer[2079] = 16'h4530;
 buffer[2080] = 16'h710F;
 buffer[2081] = 16'h1036;
 buffer[2082] = 16'h6106;
 buffer[2083] = 16'h6F62;
 buffer[2084] = 16'h7472;
 buffer[2085] = 16'h0031;
 buffer[2086] = 16'h4501;
 buffer[2087] = 16'h4542;
 buffer[2088] = 16'h803F;
 buffer[2089] = 16'h44C7;
 buffer[2090] = 16'h4529;
 buffer[2091] = 16'hFE8C;
 buffer[2092] = 16'h43BC;
 buffer[2093] = 16'h081F;
 buffer[2094] = 16'h1044;
 buffer[2095] = 16'h3C49;
 buffer[2096] = 16'h613F;
 buffer[2097] = 16'h6F62;
 buffer[2098] = 16'h7472;
 buffer[2099] = 16'h3E22;
 buffer[2100] = 16'h2837;
 buffer[2101] = 16'h4530;
 buffer[2102] = 16'h0826;
 buffer[2103] = 16'h081F;
 buffer[2104] = 16'h105E;
 buffer[2105] = 16'h6606;
 buffer[2106] = 16'h726F;
 buffer[2107] = 16'h6567;
 buffer[2108] = 16'h0074;
 buffer[2109] = 16'h474A;
 buffer[2110] = 16'h47C6;
 buffer[2111] = 16'h4264;
 buffer[2112] = 16'h284F;
 buffer[2113] = 16'h4351;
 buffer[2114] = 16'h6081;
 buffer[2115] = 16'hFEAC;
 buffer[2116] = 16'h6023;
 buffer[2117] = 16'h6103;
 buffer[2118] = 16'h6C00;
 buffer[2119] = 16'h6081;
 buffer[2120] = 16'hFE90;
 buffer[2121] = 16'h6023;
 buffer[2122] = 16'h6103;
 buffer[2123] = 16'hFEAE;
 buffer[2124] = 16'h6023;
 buffer[2125] = 16'h6103;
 buffer[2126] = 16'h710F;
 buffer[2127] = 16'h0826;
 buffer[2128] = 16'h1072;
 buffer[2129] = 16'h240A;
 buffer[2130] = 16'h6E69;
 buffer[2131] = 16'h6574;
 buffer[2132] = 16'h7072;
 buffer[2133] = 16'h6572;
 buffer[2134] = 16'h0074;
 buffer[2135] = 16'h47C6;
 buffer[2136] = 16'h4264;
 buffer[2137] = 16'h2867;
 buffer[2138] = 16'h6C00;
 buffer[2139] = 16'h8040;
 buffer[2140] = 16'h6303;
 buffer[2141] = 16'h4834;
 buffer[2142] = 16'h630C;
 buffer[2143] = 16'h6D6F;
 buffer[2144] = 16'h6970;
 buffer[2145] = 16'h656C;
 buffer[2146] = 16'h6F2D;
 buffer[2147] = 16'h6C6E;
 buffer[2148] = 16'h0079;
 buffer[2149] = 16'h0172;
 buffer[2150] = 16'h086B;
 buffer[2151] = 16'h445F;
 buffer[2152] = 16'h286A;
 buffer[2153] = 16'h700C;
 buffer[2154] = 16'h0826;
 buffer[2155] = 16'h10A2;
 buffer[2156] = 16'h5B81;
 buffer[2157] = 16'h90AE;
 buffer[2158] = 16'hFE8A;
 buffer[2159] = 16'h6023;
 buffer[2160] = 16'h710F;
 buffer[2161] = 16'h10D8;
 buffer[2162] = 16'h2E03;
 buffer[2163] = 16'h6B6F;
 buffer[2164] = 16'h90AE;
 buffer[2165] = 16'hFE8A;
 buffer[2166] = 16'h6C00;
 buffer[2167] = 16'h6703;
 buffer[2168] = 16'h287C;
 buffer[2169] = 16'h4547;
 buffer[2170] = 16'h2003;
 buffer[2171] = 16'h6B6F;
 buffer[2172] = 16'h0529;
 buffer[2173] = 16'h10E4;
 buffer[2174] = 16'h6504;
 buffer[2175] = 16'h6176;
 buffer[2176] = 16'h006C;
 buffer[2177] = 16'h474A;
 buffer[2178] = 16'h6081;
 buffer[2179] = 16'h417E;
 buffer[2180] = 16'h2888;
 buffer[2181] = 16'hFE8A;
 buffer[2182] = 16'h43BC;
 buffer[2183] = 16'h0881;
 buffer[2184] = 16'h6103;
 buffer[2185] = 16'h0874;
 buffer[2186] = 16'h10FC;
 buffer[2187] = 16'h2445;
 buffer[2188] = 16'h7665;
 buffer[2189] = 16'h6C61;
 buffer[2190] = 16'hFE84;
 buffer[2191] = 16'h6C00;
 buffer[2192] = 16'h6147;
 buffer[2193] = 16'hFE86;
 buffer[2194] = 16'h6C00;
 buffer[2195] = 16'h6147;
 buffer[2196] = 16'hFE88;
 buffer[2197] = 16'h6C00;
 buffer[2198] = 16'h6147;
 buffer[2199] = 16'hFE84;
 buffer[2200] = 16'h8000;
 buffer[2201] = 16'h6180;
 buffer[2202] = 16'h6023;
 buffer[2203] = 16'h6103;
 buffer[2204] = 16'hFE86;
 buffer[2205] = 16'h6023;
 buffer[2206] = 16'h6103;
 buffer[2207] = 16'hFE88;
 buffer[2208] = 16'h6023;
 buffer[2209] = 16'h6103;
 buffer[2210] = 16'h4881;
 buffer[2211] = 16'h6B8D;
 buffer[2212] = 16'hFE88;
 buffer[2213] = 16'h6023;
 buffer[2214] = 16'h6103;
 buffer[2215] = 16'h6B8D;
 buffer[2216] = 16'hFE86;
 buffer[2217] = 16'h6023;
 buffer[2218] = 16'h6103;
 buffer[2219] = 16'h6B8D;
 buffer[2220] = 16'hFE84;
 buffer[2221] = 16'h6023;
 buffer[2222] = 16'h710F;
 buffer[2223] = 16'h1116;
 buffer[2224] = 16'h7006;
 buffer[2225] = 16'h6572;
 buffer[2226] = 16'h6573;
 buffer[2227] = 16'h0074;
 buffer[2228] = 16'hFF00;
 buffer[2229] = 16'hFE86;
 buffer[2230] = 16'h434B;
 buffer[2231] = 16'h6023;
 buffer[2232] = 16'h710F;
 buffer[2233] = 16'h1160;
 buffer[2234] = 16'h7104;
 buffer[2235] = 16'h6975;
 buffer[2236] = 16'h0074;
 buffer[2237] = 16'h486D;
 buffer[2238] = 16'h480E;
 buffer[2239] = 16'h4881;
 buffer[2240] = 16'h08BE;
 buffer[2241] = 16'h700C;
 buffer[2242] = 16'h1174;
 buffer[2243] = 16'h6105;
 buffer[2244] = 16'h6F62;
 buffer[2245] = 16'h7472;
 buffer[2246] = 16'h6103;
 buffer[2247] = 16'h48B4;
 buffer[2248] = 16'h4874;
 buffer[2249] = 16'h08BD;
 buffer[2250] = 16'h1186;
 buffer[2251] = 16'h2701;
 buffer[2252] = 16'h474A;
 buffer[2253] = 16'h47C6;
 buffer[2254] = 16'h28D0;
 buffer[2255] = 16'h700C;
 buffer[2256] = 16'h0826;
 buffer[2257] = 16'h1196;
 buffer[2258] = 16'h6105;
 buffer[2259] = 16'h6C6C;
 buffer[2260] = 16'h746F;
 buffer[2261] = 16'h439B;
 buffer[2262] = 16'hFEAC;
 buffer[2263] = 16'h0370;
 buffer[2264] = 16'h11A4;
 buffer[2265] = 16'h2C01;
 buffer[2266] = 16'h4394;
 buffer[2267] = 16'h6081;
 buffer[2268] = 16'h434B;
 buffer[2269] = 16'hFEAC;
 buffer[2270] = 16'h6023;
 buffer[2271] = 16'h6103;
 buffer[2272] = 16'h6023;
 buffer[2273] = 16'h710F;
 buffer[2274] = 16'h11B2;
 buffer[2275] = 16'h6345;
 buffer[2276] = 16'h6C61;
 buffer[2277] = 16'h2C6C;
 buffer[2278] = 16'h8001;
 buffer[2279] = 16'h6903;
 buffer[2280] = 16'hC000;
 buffer[2281] = 16'h6403;
 buffer[2282] = 16'h08DA;
 buffer[2283] = 16'h11C6;
 buffer[2284] = 16'h3F47;
 buffer[2285] = 16'h7262;
 buffer[2286] = 16'h6E61;
 buffer[2287] = 16'h6863;
 buffer[2288] = 16'h8001;
 buffer[2289] = 16'h6903;
 buffer[2290] = 16'hA000;
 buffer[2291] = 16'h6403;
 buffer[2292] = 16'h08DA;
 buffer[2293] = 16'h11D8;
 buffer[2294] = 16'h6246;
 buffer[2295] = 16'h6172;
 buffer[2296] = 16'h636E;
 buffer[2297] = 16'h0068;
 buffer[2298] = 16'h8001;
 buffer[2299] = 16'h6903;
 buffer[2300] = 16'h8000;
 buffer[2301] = 16'h6403;
 buffer[2302] = 16'h08DA;
 buffer[2303] = 16'h11EC;
 buffer[2304] = 16'h5B89;
 buffer[2305] = 16'h6F63;
 buffer[2306] = 16'h706D;
 buffer[2307] = 16'h6C69;
 buffer[2308] = 16'h5D65;
 buffer[2309] = 16'h48CC;
 buffer[2310] = 16'h08E6;
 buffer[2311] = 16'h1200;
 buffer[2312] = 16'h6347;
 buffer[2313] = 16'h6D6F;
 buffer[2314] = 16'h6970;
 buffer[2315] = 16'h656C;
 buffer[2316] = 16'h6B8D;
 buffer[2317] = 16'h6081;
 buffer[2318] = 16'h6C00;
 buffer[2319] = 16'h48DA;
 buffer[2320] = 16'h434B;
 buffer[2321] = 16'h6147;
 buffer[2322] = 16'h700C;
 buffer[2323] = 16'h1210;
 buffer[2324] = 16'h7287;
 buffer[2325] = 16'h6365;
 buffer[2326] = 16'h7275;
 buffer[2327] = 16'h6573;
 buffer[2328] = 16'hFEAE;
 buffer[2329] = 16'h6C00;
 buffer[2330] = 16'h4750;
 buffer[2331] = 16'h08E6;
 buffer[2332] = 16'h1228;
 buffer[2333] = 16'h7004;
 buffer[2334] = 16'h6369;
 buffer[2335] = 16'h006B;
 buffer[2336] = 16'h6081;
 buffer[2337] = 16'h6410;
 buffer[2338] = 16'h6410;
 buffer[2339] = 16'h80C0;
 buffer[2340] = 16'h6203;
 buffer[2341] = 16'h6147;
 buffer[2342] = 16'h700C;
 buffer[2343] = 16'h123A;
 buffer[2344] = 16'h6C87;
 buffer[2345] = 16'h7469;
 buffer[2346] = 16'h7265;
 buffer[2347] = 16'h6C61;
 buffer[2348] = 16'h6081;
 buffer[2349] = 16'hFFFF;
 buffer[2350] = 16'h6600;
 buffer[2351] = 16'h6303;
 buffer[2352] = 16'h2938;
 buffer[2353] = 16'h8000;
 buffer[2354] = 16'h6600;
 buffer[2355] = 16'h6503;
 buffer[2356] = 16'h492C;
 buffer[2357] = 16'h490C;
 buffer[2358] = 16'h6600;
 buffer[2359] = 16'h093C;
 buffer[2360] = 16'hFFFF;
 buffer[2361] = 16'h6600;
 buffer[2362] = 16'h6403;
 buffer[2363] = 16'h08DA;
 buffer[2364] = 16'h700C;
 buffer[2365] = 16'h1250;
 buffer[2366] = 16'h5B83;
 buffer[2367] = 16'h5D27;
 buffer[2368] = 16'h48CC;
 buffer[2369] = 16'h092C;
 buffer[2370] = 16'h127C;
 buffer[2371] = 16'h2403;
 buffer[2372] = 16'h222C;
 buffer[2373] = 16'h8022;
 buffer[2374] = 16'h4718;
 buffer[2375] = 16'h4394;
 buffer[2376] = 16'h45CE;
 buffer[2377] = 16'h438C;
 buffer[2378] = 16'h6203;
 buffer[2379] = 16'h439B;
 buffer[2380] = 16'hFEAC;
 buffer[2381] = 16'h6023;
 buffer[2382] = 16'h710F;
 buffer[2383] = 16'h1286;
 buffer[2384] = 16'h66C3;
 buffer[2385] = 16'h726F;
 buffer[2386] = 16'h490C;
 buffer[2387] = 16'h4112;
 buffer[2388] = 16'h0394;
 buffer[2389] = 16'h12A0;
 buffer[2390] = 16'h62C5;
 buffer[2391] = 16'h6765;
 buffer[2392] = 16'h6E69;
 buffer[2393] = 16'h0394;
 buffer[2394] = 16'h12AC;
 buffer[2395] = 16'h2846;
 buffer[2396] = 16'h656E;
 buffer[2397] = 16'h7478;
 buffer[2398] = 16'h0029;
 buffer[2399] = 16'h6B8D;
 buffer[2400] = 16'h6B8D;
 buffer[2401] = 16'h4264;
 buffer[2402] = 16'h2968;
 buffer[2403] = 16'h6A00;
 buffer[2404] = 16'h6147;
 buffer[2405] = 16'h6C00;
 buffer[2406] = 16'h6147;
 buffer[2407] = 16'h700C;
 buffer[2408] = 16'h434B;
 buffer[2409] = 16'h6147;
 buffer[2410] = 16'h700C;
 buffer[2411] = 16'h12B6;
 buffer[2412] = 16'h6EC4;
 buffer[2413] = 16'h7865;
 buffer[2414] = 16'h0074;
 buffer[2415] = 16'h490C;
 buffer[2416] = 16'h495F;
 buffer[2417] = 16'h08DA;
 buffer[2418] = 16'h12D8;
 buffer[2419] = 16'h2844;
 buffer[2420] = 16'h6F64;
 buffer[2421] = 16'h0029;
 buffer[2422] = 16'h6B8D;
 buffer[2423] = 16'h6081;
 buffer[2424] = 16'h6147;
 buffer[2425] = 16'h6180;
 buffer[2426] = 16'h426B;
 buffer[2427] = 16'h6147;
 buffer[2428] = 16'h6147;
 buffer[2429] = 16'h434B;
 buffer[2430] = 16'h6147;
 buffer[2431] = 16'h700C;
 buffer[2432] = 16'h12E6;
 buffer[2433] = 16'h64C2;
 buffer[2434] = 16'h006F;
 buffer[2435] = 16'h490C;
 buffer[2436] = 16'h4976;
 buffer[2437] = 16'h8000;
 buffer[2438] = 16'h48DA;
 buffer[2439] = 16'h0394;
 buffer[2440] = 16'h1302;
 buffer[2441] = 16'h2847;
 buffer[2442] = 16'h656C;
 buffer[2443] = 16'h7661;
 buffer[2444] = 16'h2965;
 buffer[2445] = 16'h6B8D;
 buffer[2446] = 16'h6103;
 buffer[2447] = 16'h6B8D;
 buffer[2448] = 16'h6103;
 buffer[2449] = 16'h6B8D;
 buffer[2450] = 16'h710F;
 buffer[2451] = 16'h1312;
 buffer[2452] = 16'h6CC5;
 buffer[2453] = 16'h6165;
 buffer[2454] = 16'h6576;
 buffer[2455] = 16'h490C;
 buffer[2456] = 16'h498D;
 buffer[2457] = 16'h700C;
 buffer[2458] = 16'h1328;
 buffer[2459] = 16'h2846;
 buffer[2460] = 16'h6F6C;
 buffer[2461] = 16'h706F;
 buffer[2462] = 16'h0029;
 buffer[2463] = 16'h6B8D;
 buffer[2464] = 16'h6B8D;
 buffer[2465] = 16'h6310;
 buffer[2466] = 16'h6B8D;
 buffer[2467] = 16'h4279;
 buffer[2468] = 16'h6213;
 buffer[2469] = 16'h29AB;
 buffer[2470] = 16'h6147;
 buffer[2471] = 16'h6147;
 buffer[2472] = 16'h6C00;
 buffer[2473] = 16'h6147;
 buffer[2474] = 16'h700C;
 buffer[2475] = 16'h6147;
 buffer[2476] = 16'h6A00;
 buffer[2477] = 16'h6147;
 buffer[2478] = 16'h434B;
 buffer[2479] = 16'h6147;
 buffer[2480] = 16'h700C;
 buffer[2481] = 16'h1336;
 buffer[2482] = 16'h2848;
 buffer[2483] = 16'h6E75;
 buffer[2484] = 16'h6F6C;
 buffer[2485] = 16'h706F;
 buffer[2486] = 16'h0029;
 buffer[2487] = 16'h6B8D;
 buffer[2488] = 16'h6B8D;
 buffer[2489] = 16'h6103;
 buffer[2490] = 16'h6B8D;
 buffer[2491] = 16'h6103;
 buffer[2492] = 16'h6B8D;
 buffer[2493] = 16'h6103;
 buffer[2494] = 16'h6147;
 buffer[2495] = 16'h700C;
 buffer[2496] = 16'h1364;
 buffer[2497] = 16'h75C6;
 buffer[2498] = 16'h6C6E;
 buffer[2499] = 16'h6F6F;
 buffer[2500] = 16'h0070;
 buffer[2501] = 16'h490C;
 buffer[2502] = 16'h49B7;
 buffer[2503] = 16'h700C;
 buffer[2504] = 16'h1382;
 buffer[2505] = 16'h2845;
 buffer[2506] = 16'h643F;
 buffer[2507] = 16'h296F;
 buffer[2508] = 16'h4279;
 buffer[2509] = 16'h6213;
 buffer[2510] = 16'h29D9;
 buffer[2511] = 16'h6B8D;
 buffer[2512] = 16'h6081;
 buffer[2513] = 16'h6147;
 buffer[2514] = 16'h6180;
 buffer[2515] = 16'h426B;
 buffer[2516] = 16'h6147;
 buffer[2517] = 16'h6147;
 buffer[2518] = 16'h434B;
 buffer[2519] = 16'h6147;
 buffer[2520] = 16'h700C;
 buffer[2521] = 16'h0273;
 buffer[2522] = 16'h700C;
 buffer[2523] = 16'h1392;
 buffer[2524] = 16'h3FC3;
 buffer[2525] = 16'h6F64;
 buffer[2526] = 16'h490C;
 buffer[2527] = 16'h49CC;
 buffer[2528] = 16'h8000;
 buffer[2529] = 16'h48DA;
 buffer[2530] = 16'h0394;
 buffer[2531] = 16'h13B8;
 buffer[2532] = 16'h6CC4;
 buffer[2533] = 16'h6F6F;
 buffer[2534] = 16'h0070;
 buffer[2535] = 16'h490C;
 buffer[2536] = 16'h499F;
 buffer[2537] = 16'h6081;
 buffer[2538] = 16'h48DA;
 buffer[2539] = 16'h490C;
 buffer[2540] = 16'h49B7;
 buffer[2541] = 16'h4351;
 buffer[2542] = 16'h4394;
 buffer[2543] = 16'h8001;
 buffer[2544] = 16'h6903;
 buffer[2545] = 16'h6180;
 buffer[2546] = 16'h6023;
 buffer[2547] = 16'h710F;
 buffer[2548] = 16'h13C8;
 buffer[2549] = 16'h2847;
 buffer[2550] = 16'h6C2B;
 buffer[2551] = 16'h6F6F;
 buffer[2552] = 16'h2970;
 buffer[2553] = 16'h6B8D;
 buffer[2554] = 16'h6180;
 buffer[2555] = 16'h6B8D;
 buffer[2556] = 16'h6B8D;
 buffer[2557] = 16'h4279;
 buffer[2558] = 16'h428F;
 buffer[2559] = 16'h6147;
 buffer[2560] = 16'h8002;
 buffer[2561] = 16'h4920;
 buffer[2562] = 16'h6B81;
 buffer[2563] = 16'h6203;
 buffer[2564] = 16'h6B81;
 buffer[2565] = 16'h6503;
 buffer[2566] = 16'h6810;
 buffer[2567] = 16'h6010;
 buffer[2568] = 16'h8003;
 buffer[2569] = 16'h4920;
 buffer[2570] = 16'h6B8D;
 buffer[2571] = 16'h6503;
 buffer[2572] = 16'h6810;
 buffer[2573] = 16'h6010;
 buffer[2574] = 16'h6403;
 buffer[2575] = 16'h2A16;
 buffer[2576] = 16'h6147;
 buffer[2577] = 16'h6203;
 buffer[2578] = 16'h6147;
 buffer[2579] = 16'h6C00;
 buffer[2580] = 16'h6147;
 buffer[2581] = 16'h700C;
 buffer[2582] = 16'h6147;
 buffer[2583] = 16'h6147;
 buffer[2584] = 16'h6103;
 buffer[2585] = 16'h434B;
 buffer[2586] = 16'h6147;
 buffer[2587] = 16'h700C;
 buffer[2588] = 16'h13EA;
 buffer[2589] = 16'h2BC5;
 buffer[2590] = 16'h6F6C;
 buffer[2591] = 16'h706F;
 buffer[2592] = 16'h490C;
 buffer[2593] = 16'h49F9;
 buffer[2594] = 16'h6081;
 buffer[2595] = 16'h48DA;
 buffer[2596] = 16'h490C;
 buffer[2597] = 16'h49B7;
 buffer[2598] = 16'h4351;
 buffer[2599] = 16'h4394;
 buffer[2600] = 16'h8001;
 buffer[2601] = 16'h6903;
 buffer[2602] = 16'h6180;
 buffer[2603] = 16'h6023;
 buffer[2604] = 16'h710F;
 buffer[2605] = 16'h143A;
 buffer[2606] = 16'h2843;
 buffer[2607] = 16'h2969;
 buffer[2608] = 16'h6B8D;
 buffer[2609] = 16'h6B8D;
 buffer[2610] = 16'h414F;
 buffer[2611] = 16'h6147;
 buffer[2612] = 16'h6147;
 buffer[2613] = 16'h700C;
 buffer[2614] = 16'h145C;
 buffer[2615] = 16'h69C1;
 buffer[2616] = 16'h490C;
 buffer[2617] = 16'h4A30;
 buffer[2618] = 16'h700C;
 buffer[2619] = 16'h146E;
 buffer[2620] = 16'h75C5;
 buffer[2621] = 16'h746E;
 buffer[2622] = 16'h6C69;
 buffer[2623] = 16'h08F0;
 buffer[2624] = 16'h1478;
 buffer[2625] = 16'h61C5;
 buffer[2626] = 16'h6167;
 buffer[2627] = 16'h6E69;
 buffer[2628] = 16'h08FA;
 buffer[2629] = 16'h1482;
 buffer[2630] = 16'h69C2;
 buffer[2631] = 16'h0066;
 buffer[2632] = 16'h4394;
 buffer[2633] = 16'h8000;
 buffer[2634] = 16'h08F0;
 buffer[2635] = 16'h148C;
 buffer[2636] = 16'h74C4;
 buffer[2637] = 16'h6568;
 buffer[2638] = 16'h006E;
 buffer[2639] = 16'h4394;
 buffer[2640] = 16'h8001;
 buffer[2641] = 16'h6903;
 buffer[2642] = 16'h6181;
 buffer[2643] = 16'h6C00;
 buffer[2644] = 16'h6403;
 buffer[2645] = 16'h6180;
 buffer[2646] = 16'h6023;
 buffer[2647] = 16'h710F;
 buffer[2648] = 16'h1498;
 buffer[2649] = 16'h72C6;
 buffer[2650] = 16'h7065;
 buffer[2651] = 16'h6165;
 buffer[2652] = 16'h0074;
 buffer[2653] = 16'h48FA;
 buffer[2654] = 16'h0A4F;
 buffer[2655] = 16'h14B2;
 buffer[2656] = 16'h73C4;
 buffer[2657] = 16'h696B;
 buffer[2658] = 16'h0070;
 buffer[2659] = 16'h4394;
 buffer[2660] = 16'h8000;
 buffer[2661] = 16'h08FA;
 buffer[2662] = 16'h14C0;
 buffer[2663] = 16'h61C3;
 buffer[2664] = 16'h7466;
 buffer[2665] = 16'h6103;
 buffer[2666] = 16'h4A63;
 buffer[2667] = 16'h4959;
 buffer[2668] = 16'h718C;
 buffer[2669] = 16'h14CE;
 buffer[2670] = 16'h65C4;
 buffer[2671] = 16'h736C;
 buffer[2672] = 16'h0065;
 buffer[2673] = 16'h4A63;
 buffer[2674] = 16'h6180;
 buffer[2675] = 16'h0A4F;
 buffer[2676] = 16'h14DC;
 buffer[2677] = 16'h77C5;
 buffer[2678] = 16'h6968;
 buffer[2679] = 16'h656C;
 buffer[2680] = 16'h4A48;
 buffer[2681] = 16'h718C;
 buffer[2682] = 16'h14EA;
 buffer[2683] = 16'h2846;
 buffer[2684] = 16'h6163;
 buffer[2685] = 16'h6573;
 buffer[2686] = 16'h0029;
 buffer[2687] = 16'h6B8D;
 buffer[2688] = 16'h6180;
 buffer[2689] = 16'h6147;
 buffer[2690] = 16'h6147;
 buffer[2691] = 16'h700C;
 buffer[2692] = 16'h14F6;
 buffer[2693] = 16'h63C4;
 buffer[2694] = 16'h7361;
 buffer[2695] = 16'h0065;
 buffer[2696] = 16'h490C;
 buffer[2697] = 16'h4A7F;
 buffer[2698] = 16'h8030;
 buffer[2699] = 16'h700C;
 buffer[2700] = 16'h150A;
 buffer[2701] = 16'h2844;
 buffer[2702] = 16'h666F;
 buffer[2703] = 16'h0029;
 buffer[2704] = 16'h6B8D;
 buffer[2705] = 16'h6B81;
 buffer[2706] = 16'h6180;
 buffer[2707] = 16'h6147;
 buffer[2708] = 16'h770F;
 buffer[2709] = 16'h151A;
 buffer[2710] = 16'h6FC2;
 buffer[2711] = 16'h0066;
 buffer[2712] = 16'h490C;
 buffer[2713] = 16'h4A90;
 buffer[2714] = 16'h0A48;
 buffer[2715] = 16'h152C;
 buffer[2716] = 16'h65C5;
 buffer[2717] = 16'h646E;
 buffer[2718] = 16'h666F;
 buffer[2719] = 16'h4A71;
 buffer[2720] = 16'h8031;
 buffer[2721] = 16'h700C;
 buffer[2722] = 16'h1538;
 buffer[2723] = 16'h2809;
 buffer[2724] = 16'h6E65;
 buffer[2725] = 16'h6364;
 buffer[2726] = 16'h7361;
 buffer[2727] = 16'h2965;
 buffer[2728] = 16'h6B8D;
 buffer[2729] = 16'h6B8D;
 buffer[2730] = 16'h6103;
 buffer[2731] = 16'h6147;
 buffer[2732] = 16'h700C;
 buffer[2733] = 16'h1546;
 buffer[2734] = 16'h65C7;
 buffer[2735] = 16'h646E;
 buffer[2736] = 16'h6163;
 buffer[2737] = 16'h6573;
 buffer[2738] = 16'h6081;
 buffer[2739] = 16'h8031;
 buffer[2740] = 16'h6703;
 buffer[2741] = 16'h2AB9;
 buffer[2742] = 16'h6103;
 buffer[2743] = 16'h4A4F;
 buffer[2744] = 16'h0AB2;
 buffer[2745] = 16'h8030;
 buffer[2746] = 16'h6213;
 buffer[2747] = 16'h4834;
 buffer[2748] = 16'h6213;
 buffer[2749] = 16'h6461;
 buffer[2750] = 16'h6320;
 buffer[2751] = 16'h7361;
 buffer[2752] = 16'h2065;
 buffer[2753] = 16'h6F63;
 buffer[2754] = 16'h736E;
 buffer[2755] = 16'h7274;
 buffer[2756] = 16'h6375;
 buffer[2757] = 16'h2E74;
 buffer[2758] = 16'h490C;
 buffer[2759] = 16'h4AA8;
 buffer[2760] = 16'h700C;
 buffer[2761] = 16'h155C;
 buffer[2762] = 16'h24C2;
 buffer[2763] = 16'h0022;
 buffer[2764] = 16'h490C;
 buffer[2765] = 16'h453D;
 buffer[2766] = 16'h0945;
 buffer[2767] = 16'h1594;
 buffer[2768] = 16'h2EC2;
 buffer[2769] = 16'h0022;
 buffer[2770] = 16'h490C;
 buffer[2771] = 16'h4547;
 buffer[2772] = 16'h0945;
 buffer[2773] = 16'h15A0;
 buffer[2774] = 16'h3E05;
 buffer[2775] = 16'h6F62;
 buffer[2776] = 16'h7964;
 buffer[2777] = 16'h034B;
 buffer[2778] = 16'h15AC;
 buffer[2779] = 16'h2844;
 buffer[2780] = 16'h6F74;
 buffer[2781] = 16'h0029;
 buffer[2782] = 16'h6B8D;
 buffer[2783] = 16'h6081;
 buffer[2784] = 16'h434B;
 buffer[2785] = 16'h6147;
 buffer[2786] = 16'h6C00;
 buffer[2787] = 16'h6023;
 buffer[2788] = 16'h710F;
 buffer[2789] = 16'h15B6;
 buffer[2790] = 16'h74C2;
 buffer[2791] = 16'h006F;
 buffer[2792] = 16'h490C;
 buffer[2793] = 16'h4ADE;
 buffer[2794] = 16'h48CC;
 buffer[2795] = 16'h4AD9;
 buffer[2796] = 16'h08DA;
 buffer[2797] = 16'h15CC;
 buffer[2798] = 16'h2845;
 buffer[2799] = 16'h742B;
 buffer[2800] = 16'h296F;
 buffer[2801] = 16'h6B8D;
 buffer[2802] = 16'h6081;
 buffer[2803] = 16'h434B;
 buffer[2804] = 16'h6147;
 buffer[2805] = 16'h6C00;
 buffer[2806] = 16'h0370;
 buffer[2807] = 16'h15DC;
 buffer[2808] = 16'h2BC3;
 buffer[2809] = 16'h6F74;
 buffer[2810] = 16'h490C;
 buffer[2811] = 16'h4AF1;
 buffer[2812] = 16'h48CC;
 buffer[2813] = 16'h4AD9;
 buffer[2814] = 16'h08DA;
 buffer[2815] = 16'h15F0;
 buffer[2816] = 16'h670B;
 buffer[2817] = 16'h7465;
 buffer[2818] = 16'h632D;
 buffer[2819] = 16'h7275;
 buffer[2820] = 16'h6572;
 buffer[2821] = 16'h746E;
 buffer[2822] = 16'hFEA8;
 buffer[2823] = 16'h7C0C;
 buffer[2824] = 16'h1600;
 buffer[2825] = 16'h730B;
 buffer[2826] = 16'h7465;
 buffer[2827] = 16'h632D;
 buffer[2828] = 16'h7275;
 buffer[2829] = 16'h6572;
 buffer[2830] = 16'h746E;
 buffer[2831] = 16'hFEA8;
 buffer[2832] = 16'h6023;
 buffer[2833] = 16'h710F;
 buffer[2834] = 16'h1612;
 buffer[2835] = 16'h640B;
 buffer[2836] = 16'h6665;
 buffer[2837] = 16'h6E69;
 buffer[2838] = 16'h7469;
 buffer[2839] = 16'h6F69;
 buffer[2840] = 16'h736E;
 buffer[2841] = 16'hFE90;
 buffer[2842] = 16'h6C00;
 buffer[2843] = 16'h0B0F;
 buffer[2844] = 16'h1626;
 buffer[2845] = 16'h3F07;
 buffer[2846] = 16'h6E75;
 buffer[2847] = 16'h7169;
 buffer[2848] = 16'h6575;
 buffer[2849] = 16'h6081;
 buffer[2850] = 16'h4B06;
 buffer[2851] = 16'h4777;
 buffer[2852] = 16'h2B2C;
 buffer[2853] = 16'h4547;
 buffer[2854] = 16'h2007;
 buffer[2855] = 16'h6572;
 buffer[2856] = 16'h6564;
 buffer[2857] = 16'h2066;
 buffer[2858] = 16'h6181;
 buffer[2859] = 16'h4542;
 buffer[2860] = 16'h710F;
 buffer[2861] = 16'h163A;
 buffer[2862] = 16'h3C05;
 buffer[2863] = 16'h2C24;
 buffer[2864] = 16'h3E6E;
 buffer[2865] = 16'h6081;
 buffer[2866] = 16'h417E;
 buffer[2867] = 16'h2B46;
 buffer[2868] = 16'h4B21;
 buffer[2869] = 16'h6081;
 buffer[2870] = 16'h438C;
 buffer[2871] = 16'h6203;
 buffer[2872] = 16'h439B;
 buffer[2873] = 16'hFEAC;
 buffer[2874] = 16'h6023;
 buffer[2875] = 16'h6103;
 buffer[2876] = 16'h6081;
 buffer[2877] = 16'hFEAE;
 buffer[2878] = 16'h6023;
 buffer[2879] = 16'h6103;
 buffer[2880] = 16'h4351;
 buffer[2881] = 16'h4B06;
 buffer[2882] = 16'h6C00;
 buffer[2883] = 16'h6180;
 buffer[2884] = 16'h6023;
 buffer[2885] = 16'h710F;
 buffer[2886] = 16'h6103;
 buffer[2887] = 16'h453D;
 buffer[2888] = 16'h6E04;
 buffer[2889] = 16'h6D61;
 buffer[2890] = 16'h0065;
 buffer[2891] = 16'h0826;
 buffer[2892] = 16'h165C;
 buffer[2893] = 16'h2403;
 buffer[2894] = 16'h6E2C;
 buffer[2895] = 16'hFEBA;
 buffer[2896] = 16'h03BC;
 buffer[2897] = 16'h169A;
 buffer[2898] = 16'h2408;
 buffer[2899] = 16'h6F63;
 buffer[2900] = 16'h706D;
 buffer[2901] = 16'h6C69;
 buffer[2902] = 16'h0065;
 buffer[2903] = 16'h47C6;
 buffer[2904] = 16'h4264;
 buffer[2905] = 16'h2B61;
 buffer[2906] = 16'h6C00;
 buffer[2907] = 16'h8080;
 buffer[2908] = 16'h6303;
 buffer[2909] = 16'h2B60;
 buffer[2910] = 16'h0172;
 buffer[2911] = 16'h0B61;
 buffer[2912] = 16'h08E6;
 buffer[2913] = 16'h445F;
 buffer[2914] = 16'h2B64;
 buffer[2915] = 16'h092C;
 buffer[2916] = 16'h0826;
 buffer[2917] = 16'h16A4;
 buffer[2918] = 16'h6186;
 buffer[2919] = 16'h6F62;
 buffer[2920] = 16'h7472;
 buffer[2921] = 16'h0022;
 buffer[2922] = 16'h490C;
 buffer[2923] = 16'h4834;
 buffer[2924] = 16'h0945;
 buffer[2925] = 16'h16CC;
 buffer[2926] = 16'h3C07;
 buffer[2927] = 16'h766F;
 buffer[2928] = 16'h7265;
 buffer[2929] = 16'h3E74;
 buffer[2930] = 16'hFEAE;
 buffer[2931] = 16'h6C00;
 buffer[2932] = 16'h4B06;
 buffer[2933] = 16'h6023;
 buffer[2934] = 16'h710F;
 buffer[2935] = 16'h16DC;
 buffer[2936] = 16'h6F05;
 buffer[2937] = 16'h6576;
 buffer[2938] = 16'h7472;
 buffer[2939] = 16'hFEBC;
 buffer[2940] = 16'h03BC;
 buffer[2941] = 16'h16F0;
 buffer[2942] = 16'h6504;
 buffer[2943] = 16'h6978;
 buffer[2944] = 16'h0074;
 buffer[2945] = 16'h6B8D;
 buffer[2946] = 16'h710F;
 buffer[2947] = 16'h16FC;
 buffer[2948] = 16'h3CC3;
 buffer[2949] = 16'h3E3B;
 buffer[2950] = 16'h490C;
 buffer[2951] = 16'h4B81;
 buffer[2952] = 16'h486D;
 buffer[2953] = 16'h4B7B;
 buffer[2954] = 16'h8000;
 buffer[2955] = 16'h4394;
 buffer[2956] = 16'h6023;
 buffer[2957] = 16'h710F;
 buffer[2958] = 16'h1708;
 buffer[2959] = 16'h3BC1;
 buffer[2960] = 16'hFEBE;
 buffer[2961] = 16'h03BC;
 buffer[2962] = 16'h171E;
 buffer[2963] = 16'h5D01;
 buffer[2964] = 16'h96AE;
 buffer[2965] = 16'hFE8A;
 buffer[2966] = 16'h6023;
 buffer[2967] = 16'h710F;
 buffer[2968] = 16'h1726;
 buffer[2969] = 16'h3A01;
 buffer[2970] = 16'h474A;
 buffer[2971] = 16'h4B4F;
 buffer[2972] = 16'h0B94;
 buffer[2973] = 16'h1732;
 buffer[2974] = 16'h6909;
 buffer[2975] = 16'h6D6D;
 buffer[2976] = 16'h6465;
 buffer[2977] = 16'h6169;
 buffer[2978] = 16'h6574;
 buffer[2979] = 16'h8080;
 buffer[2980] = 16'hFEAE;
 buffer[2981] = 16'h6C00;
 buffer[2982] = 16'h6C00;
 buffer[2983] = 16'h6403;
 buffer[2984] = 16'hFEAE;
 buffer[2985] = 16'h6C00;
 buffer[2986] = 16'h6023;
 buffer[2987] = 16'h710F;
 buffer[2988] = 16'h173C;
 buffer[2989] = 16'h7504;
 buffer[2990] = 16'h6573;
 buffer[2991] = 16'h0072;
 buffer[2992] = 16'h474A;
 buffer[2993] = 16'h4B4F;
 buffer[2994] = 16'h4B7B;
 buffer[2995] = 16'h490C;
 buffer[2996] = 16'h41D2;
 buffer[2997] = 16'h08DA;
 buffer[2998] = 16'h175A;
 buffer[2999] = 16'h3C08;
 buffer[3000] = 16'h7263;
 buffer[3001] = 16'h6165;
 buffer[3002] = 16'h6574;
 buffer[3003] = 16'h003E;
 buffer[3004] = 16'h474A;
 buffer[3005] = 16'h4B4F;
 buffer[3006] = 16'h4B7B;
 buffer[3007] = 16'h838C;
 buffer[3008] = 16'h08E6;
 buffer[3009] = 16'h176E;
 buffer[3010] = 16'h6306;
 buffer[3011] = 16'h6572;
 buffer[3012] = 16'h7461;
 buffer[3013] = 16'h0065;
 buffer[3014] = 16'hFEC0;
 buffer[3015] = 16'h03BC;
 buffer[3016] = 16'h1784;
 buffer[3017] = 16'h7608;
 buffer[3018] = 16'h7261;
 buffer[3019] = 16'h6169;
 buffer[3020] = 16'h6C62;
 buffer[3021] = 16'h0065;
 buffer[3022] = 16'h4BC6;
 buffer[3023] = 16'h8000;
 buffer[3024] = 16'h08DA;
 buffer[3025] = 16'h1792;
 buffer[3026] = 16'h3209;
 buffer[3027] = 16'h6176;
 buffer[3028] = 16'h6972;
 buffer[3029] = 16'h6261;
 buffer[3030] = 16'h656C;
 buffer[3031] = 16'h4BC6;
 buffer[3032] = 16'h8000;
 buffer[3033] = 16'h48DA;
 buffer[3034] = 16'h8001;
 buffer[3035] = 16'h4357;
 buffer[3036] = 16'h08D5;
 buffer[3037] = 16'h17A4;
 buffer[3038] = 16'h2847;
 buffer[3039] = 16'h6F64;
 buffer[3040] = 16'h7365;
 buffer[3041] = 16'h293E;
 buffer[3042] = 16'h6B8D;
 buffer[3043] = 16'h8001;
 buffer[3044] = 16'h6903;
 buffer[3045] = 16'h4394;
 buffer[3046] = 16'h8001;
 buffer[3047] = 16'h6903;
 buffer[3048] = 16'hFEAE;
 buffer[3049] = 16'h6C00;
 buffer[3050] = 16'h4750;
 buffer[3051] = 16'h6081;
 buffer[3052] = 16'h434B;
 buffer[3053] = 16'hFFFF;
 buffer[3054] = 16'h6600;
 buffer[3055] = 16'h6403;
 buffer[3056] = 16'h48DA;
 buffer[3057] = 16'h6023;
 buffer[3058] = 16'h6103;
 buffer[3059] = 16'h08DA;
 buffer[3060] = 16'h17BC;
 buffer[3061] = 16'h630C;
 buffer[3062] = 16'h6D6F;
 buffer[3063] = 16'h6970;
 buffer[3064] = 16'h656C;
 buffer[3065] = 16'h6F2D;
 buffer[3066] = 16'h6C6E;
 buffer[3067] = 16'h0079;
 buffer[3068] = 16'h8040;
 buffer[3069] = 16'hFEAE;
 buffer[3070] = 16'h6C00;
 buffer[3071] = 16'h6C00;
 buffer[3072] = 16'h6403;
 buffer[3073] = 16'hFEAE;
 buffer[3074] = 16'h6C00;
 buffer[3075] = 16'h6023;
 buffer[3076] = 16'h710F;
 buffer[3077] = 16'h17EA;
 buffer[3078] = 16'h6485;
 buffer[3079] = 16'h656F;
 buffer[3080] = 16'h3E73;
 buffer[3081] = 16'h490C;
 buffer[3082] = 16'h4BE2;
 buffer[3083] = 16'h700C;
 buffer[3084] = 16'h180C;
 buffer[3085] = 16'h6304;
 buffer[3086] = 16'h6168;
 buffer[3087] = 16'h0072;
 buffer[3088] = 16'h435C;
 buffer[3089] = 16'h4742;
 buffer[3090] = 16'h6310;
 buffer[3091] = 16'h017E;
 buffer[3092] = 16'h181A;
 buffer[3093] = 16'h5B86;
 buffer[3094] = 16'h6863;
 buffer[3095] = 16'h7261;
 buffer[3096] = 16'h005D;
 buffer[3097] = 16'h4C10;
 buffer[3098] = 16'h092C;
 buffer[3099] = 16'h182A;
 buffer[3100] = 16'h6308;
 buffer[3101] = 16'h6E6F;
 buffer[3102] = 16'h7473;
 buffer[3103] = 16'h6E61;
 buffer[3104] = 16'h0074;
 buffer[3105] = 16'h4BC6;
 buffer[3106] = 16'h48DA;
 buffer[3107] = 16'h4BE2;
 buffer[3108] = 16'h7C0C;
 buffer[3109] = 16'h1838;
 buffer[3110] = 16'h6405;
 buffer[3111] = 16'h6665;
 buffer[3112] = 16'h7265;
 buffer[3113] = 16'h4BC6;
 buffer[3114] = 16'h8000;
 buffer[3115] = 16'h48DA;
 buffer[3116] = 16'h4BE2;
 buffer[3117] = 16'h6C00;
 buffer[3118] = 16'h4264;
 buffer[3119] = 16'h8000;
 buffer[3120] = 16'h6703;
 buffer[3121] = 16'h4834;
 buffer[3122] = 16'h750D;
 buffer[3123] = 16'h696E;
 buffer[3124] = 16'h696E;
 buffer[3125] = 16'h6974;
 buffer[3126] = 16'h6C61;
 buffer[3127] = 16'h7A69;
 buffer[3128] = 16'h6465;
 buffer[3129] = 16'h0172;
 buffer[3130] = 16'h184C;
 buffer[3131] = 16'h6982;
 buffer[3132] = 16'h0073;
 buffer[3133] = 16'h48CC;
 buffer[3134] = 16'h4AD9;
 buffer[3135] = 16'h6023;
 buffer[3136] = 16'h710F;
 buffer[3137] = 16'h1876;
 buffer[3138] = 16'h2E03;
 buffer[3139] = 16'h6469;
 buffer[3140] = 16'h4264;
 buffer[3141] = 16'h2C4A;
 buffer[3142] = 16'h438C;
 buffer[3143] = 16'h801F;
 buffer[3144] = 16'h6303;
 buffer[3145] = 16'h0519;
 buffer[3146] = 16'h4529;
 buffer[3147] = 16'h4547;
 buffer[3148] = 16'h7B08;
 buffer[3149] = 16'h6F6E;
 buffer[3150] = 16'h616E;
 buffer[3151] = 16'h656D;
 buffer[3152] = 16'h007D;
 buffer[3153] = 16'h700C;
 buffer[3154] = 16'h1884;
 buffer[3155] = 16'h7708;
 buffer[3156] = 16'h726F;
 buffer[3157] = 16'h6C64;
 buffer[3158] = 16'h7369;
 buffer[3159] = 16'h0074;
 buffer[3160] = 16'h43AA;
 buffer[3161] = 16'h4394;
 buffer[3162] = 16'h8000;
 buffer[3163] = 16'h48DA;
 buffer[3164] = 16'h6081;
 buffer[3165] = 16'hFEA8;
 buffer[3166] = 16'h434B;
 buffer[3167] = 16'h6081;
 buffer[3168] = 16'h6C00;
 buffer[3169] = 16'h48DA;
 buffer[3170] = 16'h6023;
 buffer[3171] = 16'h6103;
 buffer[3172] = 16'h8000;
 buffer[3173] = 16'h08DA;
 buffer[3174] = 16'h18A6;
 buffer[3175] = 16'h6F06;
 buffer[3176] = 16'h6472;
 buffer[3177] = 16'h7265;
 buffer[3178] = 16'h0040;
 buffer[3179] = 16'h6081;
 buffer[3180] = 16'h6C00;
 buffer[3181] = 16'h6081;
 buffer[3182] = 16'h2C75;
 buffer[3183] = 16'h6147;
 buffer[3184] = 16'h434B;
 buffer[3185] = 16'h4C6B;
 buffer[3186] = 16'h6B8D;
 buffer[3187] = 16'h6180;
 buffer[3188] = 16'h731C;
 buffer[3189] = 16'h700F;
 buffer[3190] = 16'h18CE;
 buffer[3191] = 16'h6709;
 buffer[3192] = 16'h7465;
 buffer[3193] = 16'h6F2D;
 buffer[3194] = 16'h6472;
 buffer[3195] = 16'h7265;
 buffer[3196] = 16'hFE90;
 buffer[3197] = 16'h0C6B;
 buffer[3198] = 16'h18EE;
 buffer[3199] = 16'h3E04;
 buffer[3200] = 16'h6977;
 buffer[3201] = 16'h0064;
 buffer[3202] = 16'h034B;
 buffer[3203] = 16'h18FE;
 buffer[3204] = 16'h2E04;
 buffer[3205] = 16'h6977;
 buffer[3206] = 16'h0064;
 buffer[3207] = 16'h4501;
 buffer[3208] = 16'h6081;
 buffer[3209] = 16'h4C82;
 buffer[3210] = 16'h434B;
 buffer[3211] = 16'h6C00;
 buffer[3212] = 16'h4264;
 buffer[3213] = 16'h2C90;
 buffer[3214] = 16'h4C44;
 buffer[3215] = 16'h710F;
 buffer[3216] = 16'h8000;
 buffer[3217] = 16'h0556;
 buffer[3218] = 16'h1908;
 buffer[3219] = 16'h2104;
 buffer[3220] = 16'h6977;
 buffer[3221] = 16'h0064;
 buffer[3222] = 16'h4C82;
 buffer[3223] = 16'h434B;
 buffer[3224] = 16'hFEAE;
 buffer[3225] = 16'h6C00;
 buffer[3226] = 16'h6180;
 buffer[3227] = 16'h6023;
 buffer[3228] = 16'h710F;
 buffer[3229] = 16'h1926;
 buffer[3230] = 16'h7604;
 buffer[3231] = 16'h636F;
 buffer[3232] = 16'h0073;
 buffer[3233] = 16'h4529;
 buffer[3234] = 16'h4547;
 buffer[3235] = 16'h7605;
 buffer[3236] = 16'h636F;
 buffer[3237] = 16'h3A73;
 buffer[3238] = 16'hFEA8;
 buffer[3239] = 16'h434B;
 buffer[3240] = 16'h6C00;
 buffer[3241] = 16'h4264;
 buffer[3242] = 16'h2CAF;
 buffer[3243] = 16'h6081;
 buffer[3244] = 16'h4C87;
 buffer[3245] = 16'h4C82;
 buffer[3246] = 16'h0CA8;
 buffer[3247] = 16'h700C;
 buffer[3248] = 16'h193C;
 buffer[3249] = 16'h6F05;
 buffer[3250] = 16'h6472;
 buffer[3251] = 16'h7265;
 buffer[3252] = 16'h4529;
 buffer[3253] = 16'h4547;
 buffer[3254] = 16'h7307;
 buffer[3255] = 16'h6165;
 buffer[3256] = 16'h6372;
 buffer[3257] = 16'h3A68;
 buffer[3258] = 16'h4C7C;
 buffer[3259] = 16'h4264;
 buffer[3260] = 16'h2CC1;
 buffer[3261] = 16'h6180;
 buffer[3262] = 16'h4C87;
 buffer[3263] = 16'h6A00;
 buffer[3264] = 16'h0CBB;
 buffer[3265] = 16'h4529;
 buffer[3266] = 16'h4547;
 buffer[3267] = 16'h6407;
 buffer[3268] = 16'h6665;
 buffer[3269] = 16'h6E69;
 buffer[3270] = 16'h3A65;
 buffer[3271] = 16'h4B06;
 buffer[3272] = 16'h0C87;
 buffer[3273] = 16'h1962;
 buffer[3274] = 16'h7309;
 buffer[3275] = 16'h7465;
 buffer[3276] = 16'h6F2D;
 buffer[3277] = 16'h6472;
 buffer[3278] = 16'h7265;
 buffer[3279] = 16'h6081;
 buffer[3280] = 16'h8000;
 buffer[3281] = 16'h6600;
 buffer[3282] = 16'h6703;
 buffer[3283] = 16'h2CD7;
 buffer[3284] = 16'h6103;
 buffer[3285] = 16'hFEA2;
 buffer[3286] = 16'h8001;
 buffer[3287] = 16'h8008;
 buffer[3288] = 16'h6181;
 buffer[3289] = 16'h6F03;
 buffer[3290] = 16'h4834;
 buffer[3291] = 16'h6F12;
 buffer[3292] = 16'h6576;
 buffer[3293] = 16'h2072;
 buffer[3294] = 16'h6973;
 buffer[3295] = 16'h657A;
 buffer[3296] = 16'h6F20;
 buffer[3297] = 16'h2066;
 buffer[3298] = 16'h7623;
 buffer[3299] = 16'h636F;
 buffer[3300] = 16'h0073;
 buffer[3301] = 16'hFE90;
 buffer[3302] = 16'h6180;
 buffer[3303] = 16'h6081;
 buffer[3304] = 16'h2CF2;
 buffer[3305] = 16'h6147;
 buffer[3306] = 16'h6180;
 buffer[3307] = 16'h6181;
 buffer[3308] = 16'h6023;
 buffer[3309] = 16'h6103;
 buffer[3310] = 16'h434B;
 buffer[3311] = 16'h6B8D;
 buffer[3312] = 16'h6A00;
 buffer[3313] = 16'h0CE7;
 buffer[3314] = 16'h6180;
 buffer[3315] = 16'h6023;
 buffer[3316] = 16'h710F;
 buffer[3317] = 16'h1994;
 buffer[3318] = 16'h6F04;
 buffer[3319] = 16'h6C6E;
 buffer[3320] = 16'h0079;
 buffer[3321] = 16'h8000;
 buffer[3322] = 16'h6600;
 buffer[3323] = 16'h0CCF;
 buffer[3324] = 16'h19EC;
 buffer[3325] = 16'h6104;
 buffer[3326] = 16'h736C;
 buffer[3327] = 16'h006F;
 buffer[3328] = 16'h4C7C;
 buffer[3329] = 16'h6181;
 buffer[3330] = 16'h6180;
 buffer[3331] = 16'h6310;
 buffer[3332] = 16'h0CCF;
 buffer[3333] = 16'h19FA;
 buffer[3334] = 16'h7008;
 buffer[3335] = 16'h6572;
 buffer[3336] = 16'h6976;
 buffer[3337] = 16'h756F;
 buffer[3338] = 16'h0073;
 buffer[3339] = 16'h4C7C;
 buffer[3340] = 16'h6180;
 buffer[3341] = 16'h6103;
 buffer[3342] = 16'h6A00;
 buffer[3343] = 16'h0CCF;
 buffer[3344] = 16'h1A0C;
 buffer[3345] = 16'h3E04;
 buffer[3346] = 16'h6F76;
 buffer[3347] = 16'h0063;
 buffer[3348] = 16'h4BC6;
 buffer[3349] = 16'h6081;
 buffer[3350] = 16'h48DA;
 buffer[3351] = 16'h4C96;
 buffer[3352] = 16'h4BE2;
 buffer[3353] = 16'h6C00;
 buffer[3354] = 16'h6147;
 buffer[3355] = 16'h4C7C;
 buffer[3356] = 16'h6180;
 buffer[3357] = 16'h6103;
 buffer[3358] = 16'h6B8D;
 buffer[3359] = 16'h6180;
 buffer[3360] = 16'h0CCF;
 buffer[3361] = 16'h1A22;
 buffer[3362] = 16'h7705;
 buffer[3363] = 16'h6469;
 buffer[3364] = 16'h666F;
 buffer[3365] = 16'h48CC;
 buffer[3366] = 16'h4AD9;
 buffer[3367] = 16'h7C0C;
 buffer[3368] = 16'h1A44;
 buffer[3369] = 16'h760A;
 buffer[3370] = 16'h636F;
 buffer[3371] = 16'h6261;
 buffer[3372] = 16'h6C75;
 buffer[3373] = 16'h7261;
 buffer[3374] = 16'h0079;
 buffer[3375] = 16'h4C58;
 buffer[3376] = 16'h0D14;
 buffer[3377] = 16'h1A52;
 buffer[3378] = 16'h5F05;
 buffer[3379] = 16'h7974;
 buffer[3380] = 16'h6570;
 buffer[3381] = 16'h6147;
 buffer[3382] = 16'h0D3A;
 buffer[3383] = 16'h438C;
 buffer[3384] = 16'h4362;
 buffer[3385] = 16'h44C7;
 buffer[3386] = 16'h6B81;
 buffer[3387] = 16'h2D40;
 buffer[3388] = 16'h6B8D;
 buffer[3389] = 16'h6A00;
 buffer[3390] = 16'h6147;
 buffer[3391] = 16'h0D37;
 buffer[3392] = 16'h6B8D;
 buffer[3393] = 16'h6103;
 buffer[3394] = 16'h710F;
 buffer[3395] = 16'h1A64;
 buffer[3396] = 16'h6403;
 buffer[3397] = 16'h2B6D;
 buffer[3398] = 16'h6181;
 buffer[3399] = 16'h8004;
 buffer[3400] = 16'h4556;
 buffer[3401] = 16'h4501;
 buffer[3402] = 16'h6147;
 buffer[3403] = 16'h0D4F;
 buffer[3404] = 16'h438C;
 buffer[3405] = 16'h8003;
 buffer[3406] = 16'h4556;
 buffer[3407] = 16'h6B81;
 buffer[3408] = 16'h2D55;
 buffer[3409] = 16'h6B8D;
 buffer[3410] = 16'h6A00;
 buffer[3411] = 16'h6147;
 buffer[3412] = 16'h0D4C;
 buffer[3413] = 16'h6B8D;
 buffer[3414] = 16'h710F;
 buffer[3415] = 16'h1A88;
 buffer[3416] = 16'h6404;
 buffer[3417] = 16'h6D75;
 buffer[3418] = 16'h0070;
 buffer[3419] = 16'hFE80;
 buffer[3420] = 16'h6C00;
 buffer[3421] = 16'h6147;
 buffer[3422] = 16'h4432;
 buffer[3423] = 16'h8010;
 buffer[3424] = 16'h4305;
 buffer[3425] = 16'h6147;
 buffer[3426] = 16'h4529;
 buffer[3427] = 16'h8010;
 buffer[3428] = 16'h4279;
 buffer[3429] = 16'h4D46;
 buffer[3430] = 16'h4155;
 buffer[3431] = 16'h8002;
 buffer[3432] = 16'h4508;
 buffer[3433] = 16'h4D35;
 buffer[3434] = 16'h6B81;
 buffer[3435] = 16'h2D70;
 buffer[3436] = 16'h6B8D;
 buffer[3437] = 16'h6A00;
 buffer[3438] = 16'h6147;
 buffer[3439] = 16'h0D62;
 buffer[3440] = 16'h6B8D;
 buffer[3441] = 16'h6103;
 buffer[3442] = 16'h6103;
 buffer[3443] = 16'h6B8D;
 buffer[3444] = 16'hFE80;
 buffer[3445] = 16'h6023;
 buffer[3446] = 16'h710F;
 buffer[3447] = 16'h1AB0;
 buffer[3448] = 16'h2E02;
 buffer[3449] = 16'h0073;
 buffer[3450] = 16'h4529;
 buffer[3451] = 16'h416A;
 buffer[3452] = 16'h6A00;
 buffer[3453] = 16'h800F;
 buffer[3454] = 16'h6303;
 buffer[3455] = 16'h6147;
 buffer[3456] = 16'h6B81;
 buffer[3457] = 16'h4920;
 buffer[3458] = 16'h4569;
 buffer[3459] = 16'h6B81;
 buffer[3460] = 16'h2D89;
 buffer[3461] = 16'h6B8D;
 buffer[3462] = 16'h6A00;
 buffer[3463] = 16'h6147;
 buffer[3464] = 16'h0D80;
 buffer[3465] = 16'h6B8D;
 buffer[3466] = 16'h6103;
 buffer[3467] = 16'h4547;
 buffer[3468] = 16'h3C04;
 buffer[3469] = 16'h6F74;
 buffer[3470] = 16'h0073;
 buffer[3471] = 16'h700C;
 buffer[3472] = 16'h1AF0;
 buffer[3473] = 16'h2807;
 buffer[3474] = 16'h6E3E;
 buffer[3475] = 16'h6D61;
 buffer[3476] = 16'h2965;
 buffer[3477] = 16'h6C00;
 buffer[3478] = 16'h4264;
 buffer[3479] = 16'h2D9F;
 buffer[3480] = 16'h4279;
 buffer[3481] = 16'h4750;
 buffer[3482] = 16'h6503;
 buffer[3483] = 16'h2D9E;
 buffer[3484] = 16'h4351;
 buffer[3485] = 16'h0D95;
 buffer[3486] = 16'h700F;
 buffer[3487] = 16'h6103;
 buffer[3488] = 16'h8000;
 buffer[3489] = 16'h700C;
 buffer[3490] = 16'h1B22;
 buffer[3491] = 16'h3E05;
 buffer[3492] = 16'h616E;
 buffer[3493] = 16'h656D;
 buffer[3494] = 16'h6147;
 buffer[3495] = 16'h4C7C;
 buffer[3496] = 16'h4264;
 buffer[3497] = 16'h2DC2;
 buffer[3498] = 16'h6180;
 buffer[3499] = 16'h6B81;
 buffer[3500] = 16'h6180;
 buffer[3501] = 16'h4D95;
 buffer[3502] = 16'h4264;
 buffer[3503] = 16'h2DC0;
 buffer[3504] = 16'h6147;
 buffer[3505] = 16'h6A00;
 buffer[3506] = 16'h6147;
 buffer[3507] = 16'h0DB5;
 buffer[3508] = 16'h6103;
 buffer[3509] = 16'h6B81;
 buffer[3510] = 16'h2DBB;
 buffer[3511] = 16'h6B8D;
 buffer[3512] = 16'h6A00;
 buffer[3513] = 16'h6147;
 buffer[3514] = 16'h0DB4;
 buffer[3515] = 16'h6B8D;
 buffer[3516] = 16'h6103;
 buffer[3517] = 16'h6B8D;
 buffer[3518] = 16'h6B8D;
 buffer[3519] = 16'h710F;
 buffer[3520] = 16'h6A00;
 buffer[3521] = 16'h0DA8;
 buffer[3522] = 16'h6B8D;
 buffer[3523] = 16'h6103;
 buffer[3524] = 16'h8000;
 buffer[3525] = 16'h700C;
 buffer[3526] = 16'h1B46;
 buffer[3527] = 16'h7303;
 buffer[3528] = 16'h6565;
 buffer[3529] = 16'h48CC;
 buffer[3530] = 16'h4529;
 buffer[3531] = 16'h6081;
 buffer[3532] = 16'h6C00;
 buffer[3533] = 16'h4264;
 buffer[3534] = 16'hF00C;
 buffer[3535] = 16'h6503;
 buffer[3536] = 16'h2DE2;
 buffer[3537] = 16'hBFFF;
 buffer[3538] = 16'h6303;
 buffer[3539] = 16'h8001;
 buffer[3540] = 16'h6D03;
 buffer[3541] = 16'h4DA6;
 buffer[3542] = 16'h4264;
 buffer[3543] = 16'h2DDB;
 buffer[3544] = 16'h4501;
 buffer[3545] = 16'h4C44;
 buffer[3546] = 16'h0DE0;
 buffer[3547] = 16'h6081;
 buffer[3548] = 16'h6C00;
 buffer[3549] = 16'hFFFF;
 buffer[3550] = 16'h6303;
 buffer[3551] = 16'h4562;
 buffer[3552] = 16'h434B;
 buffer[3553] = 16'h0DCB;
 buffer[3554] = 16'h0273;
 buffer[3555] = 16'h1B8E;
 buffer[3556] = 16'h2807;
 buffer[3557] = 16'h6F77;
 buffer[3558] = 16'h6472;
 buffer[3559] = 16'h2973;
 buffer[3560] = 16'h4529;
 buffer[3561] = 16'h6C00;
 buffer[3562] = 16'h4264;
 buffer[3563] = 16'h2DF1;
 buffer[3564] = 16'h6081;
 buffer[3565] = 16'h4C44;
 buffer[3566] = 16'h4501;
 buffer[3567] = 16'h4351;
 buffer[3568] = 16'h0DE9;
 buffer[3569] = 16'h700C;
 buffer[3570] = 16'h1BC8;
 buffer[3571] = 16'h7705;
 buffer[3572] = 16'h726F;
 buffer[3573] = 16'h7364;
 buffer[3574] = 16'h4C7C;
 buffer[3575] = 16'h4264;
 buffer[3576] = 16'h2E04;
 buffer[3577] = 16'h6180;
 buffer[3578] = 16'h4529;
 buffer[3579] = 16'h4529;
 buffer[3580] = 16'h4547;
 buffer[3581] = 16'h3A01;
 buffer[3582] = 16'h6081;
 buffer[3583] = 16'h4C87;
 buffer[3584] = 16'h4529;
 buffer[3585] = 16'h4DE8;
 buffer[3586] = 16'h6A00;
 buffer[3587] = 16'h0DF7;
 buffer[3588] = 16'h700C;
 buffer[3589] = 16'h1BE6;
 buffer[3590] = 16'h7603;
 buffer[3591] = 16'h7265;
 buffer[3592] = 16'h8001;
 buffer[3593] = 16'h8100;
 buffer[3594] = 16'h4329;
 buffer[3595] = 16'h8006;
 buffer[3596] = 16'h720F;
 buffer[3597] = 16'h1C0C;
 buffer[3598] = 16'h6802;
 buffer[3599] = 16'h0069;
 buffer[3600] = 16'h4529;
 buffer[3601] = 16'h4547;
 buffer[3602] = 16'h650C;
 buffer[3603] = 16'h6F66;
 buffer[3604] = 16'h7472;
 buffer[3605] = 16'h2068;
 buffer[3606] = 16'h316A;
 buffer[3607] = 16'h202B;
 buffer[3608] = 16'h0076;
 buffer[3609] = 16'hFE80;
 buffer[3610] = 16'h6C00;
 buffer[3611] = 16'h4432;
 buffer[3612] = 16'h4E08;
 buffer[3613] = 16'h43F4;
 buffer[3614] = 16'h4406;
 buffer[3615] = 16'h4406;
 buffer[3616] = 16'h802E;
 buffer[3617] = 16'h43FC;
 buffer[3618] = 16'h4406;
 buffer[3619] = 16'h441E;
 buffer[3620] = 16'h4519;
 buffer[3621] = 16'hFE80;
 buffer[3622] = 16'h6023;
 buffer[3623] = 16'h6103;
 buffer[3624] = 16'h0529;
 buffer[3625] = 16'h1C1C;
 buffer[3626] = 16'h6304;
 buffer[3627] = 16'h6C6F;
 buffer[3628] = 16'h0064;
 buffer[3629] = 16'h8002;
 buffer[3630] = 16'hFE80;
 buffer[3631] = 16'h8042;
 buffer[3632] = 16'h45B7;
 buffer[3633] = 16'h48B4;
 buffer[3634] = 16'hFEA2;
 buffer[3635] = 16'h6081;
 buffer[3636] = 16'hFE90;
 buffer[3637] = 16'h6023;
 buffer[3638] = 16'h6103;
 buffer[3639] = 16'h6081;
 buffer[3640] = 16'hFEA8;
 buffer[3641] = 16'h4379;
 buffer[3642] = 16'h4B7B;
 buffer[3643] = 16'hC000;
 buffer[3644] = 16'h434B;
 buffer[3645] = 16'h6081;
 buffer[3646] = 16'h4351;
 buffer[3647] = 16'h6C00;
 buffer[3648] = 16'h488E;
 buffer[3649] = 16'hFEB4;
 buffer[3650] = 16'h43BC;
 buffer[3651] = 16'h48BD;
 buffer[3652] = 16'h0E2D;
end

endmodule

module M_main_mem_ram(
input      [0:0]             in_ram_wenable0,
input       [15:0]     in_ram_wdata0,
input      [14:0]                in_ram_addr0,
input      [0:0]             in_ram_wenable1,
input      [15:0]                 in_ram_wdata1,
input      [14:0]                in_ram_addr1,
output reg  [15:0]     out_ram_rdata0,
output reg  [15:0]     out_ram_rdata1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[32767:0];
always @(posedge clock0) begin
  if (in_ram_wenable0) begin
    buffer[in_ram_addr0] <= in_ram_wdata0;
  end else begin
    out_ram_rdata0 <= buffer[in_ram_addr0];
  end
end
always @(posedge clock1) begin
  if (in_ram_wenable1) begin
    buffer[in_ram_addr1] <= in_ram_wdata1;
  end else begin
    out_ram_rdata1 <= buffer[in_ram_addr1];
  end
end

endmodule

module M_main_mem_uartInBuffer(
input      [0:0]             in_uartInBuffer_wenable0,
input       [7:0]     in_uartInBuffer_wdata0,
input      [7:0]                in_uartInBuffer_addr0,
input      [0:0]             in_uartInBuffer_wenable1,
input      [7:0]                 in_uartInBuffer_wdata1,
input      [7:0]                in_uartInBuffer_addr1,
output reg  [7:0]     out_uartInBuffer_rdata0,
output reg  [7:0]     out_uartInBuffer_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[255:0];
always @(posedge clock0) begin
  if (in_uartInBuffer_wenable0) begin
    buffer[in_uartInBuffer_addr0] <= in_uartInBuffer_wdata0;
  end else begin
    out_uartInBuffer_rdata0 <= buffer[in_uartInBuffer_addr0];
  end
end
always @(posedge clock1) begin
  if (in_uartInBuffer_wenable1) begin
    buffer[in_uartInBuffer_addr1] <= in_uartInBuffer_wdata1;
  end else begin
    out_uartInBuffer_rdata1 <= buffer[in_uartInBuffer_addr1];
  end
end

endmodule

module M_main_mem_uartOutBuffer(
input      [0:0]             in_uartOutBuffer_wenable0,
input       [7:0]     in_uartOutBuffer_wdata0,
input      [7:0]                in_uartOutBuffer_addr0,
input      [0:0]             in_uartOutBuffer_wenable1,
input      [7:0]                 in_uartOutBuffer_wdata1,
input      [7:0]                in_uartOutBuffer_addr1,
output reg  [7:0]     out_uartOutBuffer_rdata0,
output reg  [7:0]     out_uartOutBuffer_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[255:0];
always @(posedge clock0) begin
  if (in_uartOutBuffer_wenable0) begin
    buffer[in_uartOutBuffer_addr0] <= in_uartOutBuffer_wdata0;
  end else begin
    out_uartOutBuffer_rdata0 <= buffer[in_uartOutBuffer_addr0];
  end
end
always @(posedge clock1) begin
  if (in_uartOutBuffer_wenable1) begin
    buffer[in_uartOutBuffer_addr1] <= in_uartOutBuffer_wdata1;
  end else begin
    out_uartOutBuffer_rdata1 <= buffer[in_uartOutBuffer_addr1];
  end
end

endmodule

module M_main (
in_buttons,
in_uart_tx_busy,
in_uart_tx_done,
in_uart_rx_data,
in_uart_rx_valid,
in_timer1hz,
out_led,
out_uart_tx_data,
out_uart_tx_valid,
out_sdram_cle,
out_sdram_dqm,
out_sdram_cs,
out_sdram_we,
out_sdram_cas,
out_sdram_ras,
out_sdram_ba,
out_sdram_a,
out_sdram_clk,
out_video_r,
out_video_g,
out_video_b,
out_video_hs,
out_video_vs,
inout_sdram_dq,
in_run,
out_done,
reset,
clock
);
input  [7:0] in_buttons;
input  [0:0] in_uart_tx_busy;
input  [0:0] in_uart_tx_done;
input  [7:0] in_uart_rx_data;
input  [0:0] in_uart_rx_valid;
input  [15:0] in_timer1hz;
output  [7:0] out_led;
output  [7:0] out_uart_tx_data;
output  [0:0] out_uart_tx_valid;
output  [0:0] out_sdram_cle;
output  [0:0] out_sdram_dqm;
output  [0:0] out_sdram_cs;
output  [0:0] out_sdram_we;
output  [0:0] out_sdram_cas;
output  [0:0] out_sdram_ras;
output  [1:0] out_sdram_ba;
output  [12:0] out_sdram_a;
output  [0:0] out_sdram_clk;
output  [5:0] out_video_r;
output  [5:0] out_video_g;
output  [5:0] out_video_b;
output  [0:0] out_video_hs;
output  [0:0] out_video_vs;
inout  [7:0] inout_sdram_dq;
input in_run;
output out_done;
input reset;
input clock;
wire _w_vga_rstcond_out;
wire _w_clk_gen_outclk_0;
wire _w_clk_gen_outclk_1;
wire _w_clk_gen_locked;
wire  [0:0] _w_vga_driver_vga_hs;
wire  [0:0] _w_vga_driver_vga_vs;
wire  [0:0] _w_vga_driver_active;
wire  [0:0] _w_vga_driver_vblank;
wire  [9:0] _w_vga_driver_vga_x;
wire  [9:0] _w_vga_driver_vga_y;
wire _w_vga_driver_done;
wire  [5:0] _w_display_pix_red;
wire  [5:0] _w_display_pix_green;
wire  [5:0] _w_display_pix_blue;
wire _w_display_done;
wire  [15:0] _w_mem_dstack_rdata;
wire  [15:0] _w_mem_rstack_rdata;
wire  [15:0] _w_mem_rom_rdata;
wire  [15:0] _w_mem_ram_rdata0;
wire  [15:0] _w_mem_ram_rdata1;
wire  [7:0] _w_mem_uartInBuffer_rdata0;
wire  [7:0] _w_mem_uartInBuffer_rdata1;
wire  [7:0] _w_mem_uartOutBuffer_rdata0;
wire  [7:0] _w_mem_uartOutBuffer_rdata1;
wire  [15:0] _c_ram_wdata1;
assign _c_ram_wdata1 = 0;
wire  [7:0] _c_uartInBuffer_wdata0;
assign _c_uartInBuffer_wdata0 = 0;
wire  [7:0] _c_uartOutBuffer_wdata0;
assign _c_uartOutBuffer_wdata0 = 0;
wire  [15:0] _w_immediate;
wire  [0:0] _w_is_alu;
wire  [0:0] _w_is_call;
wire  [0:0] _w_is_lit;
wire  [0:0] _w_dstackWrite;
wire  [0:0] _w_rstackWrite;
wire  [7:0] _w_ddelta;
wire  [7:0] _w_rdelta;
wire  [12:0] _w_pcPlusOne;

reg  [15:0] _d_instruction;
reg  [15:0] _q_instruction;
reg  [12:0] _d_pc;
reg  [12:0] _q_pc;
reg  [12:0] _d_newPC;
reg  [12:0] _q_newPC;
reg  [0:0] _d_dstack_wenable;
reg  [0:0] _q_dstack_wenable;
reg  [15:0] _d_dstack_wdata;
reg  [15:0] _q_dstack_wdata;
reg  [7:0] _d_dstack_addr;
reg  [7:0] _q_dstack_addr;
reg  [15:0] _d_stackTop;
reg  [15:0] _q_stackTop;
reg  [7:0] _d_dsp;
reg  [7:0] _q_dsp;
reg  [7:0] _d_newDSP;
reg  [7:0] _q_newDSP;
reg  [15:0] _d_newStackTop;
reg  [15:0] _q_newStackTop;
reg  [0:0] _d_rstack_wenable;
reg  [0:0] _q_rstack_wenable;
reg  [15:0] _d_rstack_wdata;
reg  [15:0] _q_rstack_wdata;
reg  [7:0] _d_rstack_addr;
reg  [7:0] _q_rstack_addr;
reg  [7:0] _d_rsp;
reg  [7:0] _q_rsp;
reg  [7:0] _d_newRSP;
reg  [7:0] _q_newRSP;
reg  [15:0] _d_rstackWData;
reg  [15:0] _q_rstackWData;
reg  [15:0] _d_stackNext;
reg  [15:0] _q_stackNext;
reg  [15:0] _d_rStackTop;
reg  [15:0] _q_rStackTop;
reg  [15:0] _d_memoryInput;
reg  [15:0] _q_memoryInput;
reg  [11:0] _d_rom_addr;
reg  [11:0] _q_rom_addr;
reg  [0:0] _d_ram_wenable0;
reg  [0:0] _q_ram_wenable0;
reg  [15:0] _d_ram_wdata0;
reg  [15:0] _q_ram_wdata0;
reg  [14:0] _d_ram_addr0;
reg  [14:0] _q_ram_addr0;
reg  [0:0] _d_ram_wenable1;
reg  [0:0] _q_ram_wenable1;
reg  [14:0] _d_ram_addr1;
reg  [14:0] _q_ram_addr1;
reg  [2:0] _d_CYCLE;
reg  [2:0] _q_CYCLE;
reg  [1:0] _d_INIT;
reg  [1:0] _q_INIT;
reg  [15:0] _d_copyaddress;
reg  [15:0] _q_copyaddress;
reg  [15:0] _d_bramREAD;
reg  [15:0] _q_bramREAD;
reg  [0:0] _d_uartInBuffer_wenable0;
reg  [0:0] _q_uartInBuffer_wenable0;
reg  [7:0] _d_uartInBuffer_addr0;
reg  [7:0] _q_uartInBuffer_addr0;
reg  [0:0] _d_uartInBuffer_wenable1;
reg  [0:0] _q_uartInBuffer_wenable1;
reg  [7:0] _d_uartInBuffer_wdata1;
reg  [7:0] _q_uartInBuffer_wdata1;
reg  [7:0] _d_uartInBuffer_addr1;
reg  [7:0] _q_uartInBuffer_addr1;
reg  [7:0] _d_uartInBufferNext;
reg  [7:0] _q_uartInBufferNext;
reg  [7:0] _d_uartInBufferTop;
reg  [7:0] _q_uartInBufferTop;
reg  [0:0] _d_uartInHold;
reg  [0:0] _q_uartInHold;
reg  [0:0] _d_uartOutBuffer_wenable0;
reg  [0:0] _q_uartOutBuffer_wenable0;
reg  [7:0] _d_uartOutBuffer_addr0;
reg  [7:0] _q_uartOutBuffer_addr0;
reg  [0:0] _d_uartOutBuffer_wenable1;
reg  [0:0] _q_uartOutBuffer_wenable1;
reg  [7:0] _d_uartOutBuffer_wdata1;
reg  [7:0] _q_uartOutBuffer_wdata1;
reg  [7:0] _d_uartOutBuffer_addr1;
reg  [7:0] _q_uartOutBuffer_addr1;
reg  [7:0] _d_uartOutBufferNext;
reg  [7:0] _q_uartOutBufferNext;
reg  [7:0] _d_uartOutBufferTop;
reg  [7:0] _q_uartOutBufferTop;
reg  [7:0] _d_newuartOutBufferTop;
reg  [7:0] _q_newuartOutBufferTop;
reg  [7:0] _d_uartOutHold;
reg  [7:0] _q_uartOutHold;
reg  [7:0] _d_led,_q_led;
reg  [7:0] _d_uart_tx_data,_q_uart_tx_data;
reg  [0:0] _d_uart_tx_valid,_q_uart_tx_valid;
reg  [0:0] _d_sdram_cle,_q_sdram_cle;
reg  [0:0] _d_sdram_dqm,_q_sdram_dqm;
reg  [0:0] _d_sdram_cs,_q_sdram_cs;
reg  [0:0] _d_sdram_we,_q_sdram_we;
reg  [0:0] _d_sdram_cas,_q_sdram_cas;
reg  [0:0] _d_sdram_ras,_q_sdram_ras;
reg  [1:0] _d_sdram_ba,_q_sdram_ba;
reg  [12:0] _d_sdram_a,_q_sdram_a;
reg  [0:0] _d_sdram_clk,_q_sdram_clk;
reg  [9:0] _d_display_gpu_x,_q_display_gpu_x;
reg  [8:0] _d_display_gpu_y,_q_display_gpu_y;
reg  [7:0] _d_display_gpu_dotset,_q_display_gpu_dotset;
reg  [0:0] _d_display_gpu_write,_q_display_gpu_write;
reg  [6:0] _d_display_tpu_x,_q_display_tpu_x;
reg  [4:0] _d_display_tpu_y,_q_display_tpu_y;
reg  [7:0] _d_display_tpu_set,_q_display_tpu_set;
reg  [1:0] _d_display_tpu_write,_q_display_tpu_write;
reg  [2:0] _d_index,_q_index;
reg  _vga_driver_run;
reg  _display_run;
assign out_led = _q_led;
assign out_uart_tx_data = _q_uart_tx_data;
assign out_uart_tx_valid = _q_uart_tx_valid;
assign out_sdram_cle = _d_sdram_cle;
assign out_sdram_dqm = _d_sdram_dqm;
assign out_sdram_cs = _d_sdram_cs;
assign out_sdram_we = _d_sdram_we;
assign out_sdram_cas = _d_sdram_cas;
assign out_sdram_ras = _d_sdram_ras;
assign out_sdram_ba = _d_sdram_ba;
assign out_sdram_a = _d_sdram_a;
assign out_sdram_clk = _d_sdram_clk;
assign out_video_r = _w_display_pix_red;
assign out_video_g = _w_display_pix_green;
assign out_video_b = _w_display_pix_blue;
assign out_video_hs = _w_vga_driver_vga_hs;
assign out_video_vs = _w_vga_driver_vga_vs;
assign out_done = (_q_index == 7);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_pc <= 0;
_q_dstack_wenable <= 0;
_q_dstack_wdata <= 0;
_q_dstack_addr <= 0;
_q_stackTop <= 0;
_q_dsp <= 0;
_q_rstack_wenable <= 0;
_q_rstack_wdata <= 0;
_q_rstack_addr <= 0;
_q_rsp <= 0;
_q_rom_addr <= 0;
_q_ram_wenable0 <= 0;
_q_ram_wdata0 <= 0;
_q_ram_addr0 <= 0;
_q_ram_wenable1 <= 0;
_q_ram_addr1 <= 0;
_q_CYCLE <= 0;
_q_INIT <= 0;
_q_copyaddress <= 0;
_q_bramREAD <= 0;
_q_uartInBuffer_wenable0 <= 0;
_q_uartInBuffer_addr0 <= 0;
_q_uartInBuffer_wenable1 <= 0;
_q_uartInBuffer_wdata1 <= 0;
_q_uartInBuffer_addr1 <= 0;
_q_uartInBufferNext <= 0;
_q_uartInBufferTop <= 0;
_q_uartInHold <= 1;
_q_uartOutBuffer_wenable0 <= 0;
_q_uartOutBuffer_addr0 <= 0;
_q_uartOutBuffer_wenable1 <= 0;
_q_uartOutBuffer_wdata1 <= 0;
_q_uartOutBuffer_addr1 <= 0;
_q_uartOutBufferNext <= 0;
_q_uartOutBufferTop <= 0;
_q_newuartOutBufferTop <= 0;
_q_uartOutHold <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_instruction <= _d_instruction;
_q_pc <= _d_pc;
_q_newPC <= _d_newPC;
_q_dstack_wenable <= _d_dstack_wenable;
_q_dstack_wdata <= _d_dstack_wdata;
_q_dstack_addr <= _d_dstack_addr;
_q_stackTop <= _d_stackTop;
_q_dsp <= _d_dsp;
_q_newDSP <= _d_newDSP;
_q_newStackTop <= _d_newStackTop;
_q_rstack_wenable <= _d_rstack_wenable;
_q_rstack_wdata <= _d_rstack_wdata;
_q_rstack_addr <= _d_rstack_addr;
_q_rsp <= _d_rsp;
_q_newRSP <= _d_newRSP;
_q_rstackWData <= _d_rstackWData;
_q_stackNext <= _d_stackNext;
_q_rStackTop <= _d_rStackTop;
_q_memoryInput <= _d_memoryInput;
_q_rom_addr <= _d_rom_addr;
_q_ram_wenable0 <= _d_ram_wenable0;
_q_ram_wdata0 <= _d_ram_wdata0;
_q_ram_addr0 <= _d_ram_addr0;
_q_ram_wenable1 <= _d_ram_wenable1;
_q_ram_addr1 <= _d_ram_addr1;
_q_CYCLE <= _d_CYCLE;
_q_INIT <= _d_INIT;
_q_copyaddress <= _d_copyaddress;
_q_bramREAD <= _d_bramREAD;
_q_uartInBuffer_wenable0 <= _d_uartInBuffer_wenable0;
_q_uartInBuffer_addr0 <= _d_uartInBuffer_addr0;
_q_uartInBuffer_wenable1 <= _d_uartInBuffer_wenable1;
_q_uartInBuffer_wdata1 <= _d_uartInBuffer_wdata1;
_q_uartInBuffer_addr1 <= _d_uartInBuffer_addr1;
_q_uartInBufferNext <= _d_uartInBufferNext;
_q_uartInBufferTop <= _d_uartInBufferTop;
_q_uartInHold <= _d_uartInHold;
_q_uartOutBuffer_wenable0 <= _d_uartOutBuffer_wenable0;
_q_uartOutBuffer_addr0 <= _d_uartOutBuffer_addr0;
_q_uartOutBuffer_wenable1 <= _d_uartOutBuffer_wenable1;
_q_uartOutBuffer_wdata1 <= _d_uartOutBuffer_wdata1;
_q_uartOutBuffer_addr1 <= _d_uartOutBuffer_addr1;
_q_uartOutBufferNext <= _d_uartOutBufferNext;
_q_uartOutBufferTop <= _d_uartOutBufferTop;
_q_newuartOutBufferTop <= _d_newuartOutBufferTop;
_q_uartOutHold <= _d_uartOutHold;
_q_index <= _d_index;
  end
_q_led <= _d_led;
_q_uart_tx_data <= _d_uart_tx_data;
_q_uart_tx_valid <= _d_uart_tx_valid;
_q_sdram_cle <= _d_sdram_cle;
_q_sdram_dqm <= _d_sdram_dqm;
_q_sdram_cs <= _d_sdram_cs;
_q_sdram_we <= _d_sdram_we;
_q_sdram_cas <= _d_sdram_cas;
_q_sdram_ras <= _d_sdram_ras;
_q_sdram_ba <= _d_sdram_ba;
_q_sdram_a <= _d_sdram_a;
_q_sdram_clk <= _d_sdram_clk;
_q_display_gpu_x <= _d_display_gpu_x;
_q_display_gpu_y <= _d_display_gpu_y;
_q_display_gpu_dotset <= _d_display_gpu_dotset;
_q_display_gpu_write <= _d_display_gpu_write;
_q_display_tpu_x <= _d_display_tpu_x;
_q_display_tpu_y <= _d_display_tpu_y;
_q_display_tpu_set <= _d_display_tpu_set;
_q_display_tpu_write <= _d_display_tpu_write;
end


reset_conditioner _vga_rstcond (
.rcclk(_w_clk_gen_outclk_1),
.in(reset),
.out(_w_vga_rstcond_out)
);

de10nano_clk_100_25 _clk_gen (
.refclk(clock),
.outclk_0(_w_clk_gen_outclk_0),
.outclk_1(_w_clk_gen_outclk_1),
.locked(_w_clk_gen_locked),
.rst(reset)
);
M_vga vga_driver (
.out_vga_hs(_w_vga_driver_vga_hs),
.out_vga_vs(_w_vga_driver_vga_vs),
.out_active(_w_vga_driver_active),
.out_vblank(_w_vga_driver_vblank),
.out_vga_x(_w_vga_driver_vga_x),
.out_vga_y(_w_vga_driver_vga_y),
.out_done(_w_vga_driver_done),
.in_run(_vga_driver_run),
.reset(_w_vga_rstcond_out),
.clock(_w_clk_gen_outclk_1)
);
M_multiplex_display display (
.in_pix_x(_w_vga_driver_vga_x),
.in_pix_y(_w_vga_driver_vga_y),
.in_pix_active(_w_vga_driver_active),
.in_pix_vblank(_w_vga_driver_vblank),
.in_gpu_x(_d_display_gpu_x),
.in_gpu_y(_d_display_gpu_y),
.in_gpu_dotset(_d_display_gpu_dotset),
.in_gpu_write(_d_display_gpu_write),
.in_tpu_x(_d_display_tpu_x),
.in_tpu_y(_d_display_tpu_y),
.in_tpu_set(_d_display_tpu_set),
.in_tpu_write(_d_display_tpu_write),
.out_pix_red(_w_display_pix_red),
.out_pix_green(_w_display_pix_green),
.out_pix_blue(_w_display_pix_blue),
.out_done(_w_display_done),
.in_run(_display_run),
.reset(_w_vga_rstcond_out),
.clock(_w_clk_gen_outclk_1)
);

M_main_mem_dstack __mem__dstack(
.clock(clock),
.in_dstack_wenable(_d_dstack_wenable),
.in_dstack_wdata(_d_dstack_wdata),
.in_dstack_addr(_d_dstack_addr),
.out_dstack_rdata(_w_mem_dstack_rdata)
);
M_main_mem_rstack __mem__rstack(
.clock(clock),
.in_rstack_wenable(_d_rstack_wenable),
.in_rstack_wdata(_d_rstack_wdata),
.in_rstack_addr(_d_rstack_addr),
.out_rstack_rdata(_w_mem_rstack_rdata)
);
M_main_mem_rom __mem__rom(
.clock(clock),
.in_rom_addr(_d_rom_addr),
.out_rom_rdata(_w_mem_rom_rdata)
);
M_main_mem_ram __mem__ram(
.clock0(clock),
.clock1(clock),
.in_ram_wenable0(_d_ram_wenable0),
.in_ram_wdata0(_d_ram_wdata0),
.in_ram_addr0(_d_ram_addr0),
.in_ram_wenable1(_d_ram_wenable1),
.in_ram_wdata1(_c_ram_wdata1),
.in_ram_addr1(_d_ram_addr1),
.out_ram_rdata0(_w_mem_ram_rdata0),
.out_ram_rdata1(_w_mem_ram_rdata1)
);
M_main_mem_uartInBuffer __mem__uartInBuffer(
.clock0(clock),
.clock1(clock),
.in_uartInBuffer_wenable0(_d_uartInBuffer_wenable0),
.in_uartInBuffer_wdata0(_c_uartInBuffer_wdata0),
.in_uartInBuffer_addr0(_d_uartInBuffer_addr0),
.in_uartInBuffer_wenable1(_d_uartInBuffer_wenable1),
.in_uartInBuffer_wdata1(_d_uartInBuffer_wdata1),
.in_uartInBuffer_addr1(_d_uartInBuffer_addr1),
.out_uartInBuffer_rdata0(_w_mem_uartInBuffer_rdata0),
.out_uartInBuffer_rdata1(_w_mem_uartInBuffer_rdata1)
);
M_main_mem_uartOutBuffer __mem__uartOutBuffer(
.clock0(clock),
.clock1(clock),
.in_uartOutBuffer_wenable0(_d_uartOutBuffer_wenable0),
.in_uartOutBuffer_wdata0(_c_uartOutBuffer_wdata0),
.in_uartOutBuffer_addr0(_d_uartOutBuffer_addr0),
.in_uartOutBuffer_wenable1(_d_uartOutBuffer_wenable1),
.in_uartOutBuffer_wdata1(_d_uartOutBuffer_wdata1),
.in_uartOutBuffer_addr1(_d_uartOutBuffer_addr1),
.out_uartOutBuffer_rdata0(_w_mem_uartOutBuffer_rdata0),
.out_uartOutBuffer_rdata1(_w_mem_uartOutBuffer_rdata1)
);

assign _w_pcPlusOne = _d_pc+1;
assign _w_rdelta = {{7{_d_instruction[3+:1]}},_d_instruction[2+:1]};
assign _w_rstackWrite = (_w_is_call|(_w_is_alu&_d_instruction[6+:1]));
assign _w_dstackWrite = (_w_is_lit|(_w_is_alu&_d_instruction[7+:1]));
assign _w_ddelta = {{7{_d_instruction[1+:1]}},_d_instruction[0+:1]};
assign _w_is_call = (_d_instruction[13+:3]==3'b010);
assign _w_is_lit = _d_instruction[15+:1];
assign _w_is_alu = (_d_instruction[13+:3]==3'b011);
assign _w_immediate = (_d_instruction[0+:15]);

always @* begin
_d_instruction = _q_instruction;
_d_pc = _q_pc;
_d_newPC = _q_newPC;
_d_dstack_wenable = _q_dstack_wenable;
_d_dstack_wdata = _q_dstack_wdata;
_d_dstack_addr = _q_dstack_addr;
_d_stackTop = _q_stackTop;
_d_dsp = _q_dsp;
_d_newDSP = _q_newDSP;
_d_newStackTop = _q_newStackTop;
_d_rstack_wenable = _q_rstack_wenable;
_d_rstack_wdata = _q_rstack_wdata;
_d_rstack_addr = _q_rstack_addr;
_d_rsp = _q_rsp;
_d_newRSP = _q_newRSP;
_d_rstackWData = _q_rstackWData;
_d_stackNext = _q_stackNext;
_d_rStackTop = _q_rStackTop;
_d_memoryInput = _q_memoryInput;
_d_rom_addr = _q_rom_addr;
_d_ram_wenable0 = _q_ram_wenable0;
_d_ram_wdata0 = _q_ram_wdata0;
_d_ram_addr0 = _q_ram_addr0;
_d_ram_wenable1 = _q_ram_wenable1;
_d_ram_addr1 = _q_ram_addr1;
_d_CYCLE = _q_CYCLE;
_d_INIT = _q_INIT;
_d_copyaddress = _q_copyaddress;
_d_bramREAD = _q_bramREAD;
_d_uartInBuffer_wenable0 = _q_uartInBuffer_wenable0;
_d_uartInBuffer_addr0 = _q_uartInBuffer_addr0;
_d_uartInBuffer_wenable1 = _q_uartInBuffer_wenable1;
_d_uartInBuffer_wdata1 = _q_uartInBuffer_wdata1;
_d_uartInBuffer_addr1 = _q_uartInBuffer_addr1;
_d_uartInBufferNext = _q_uartInBufferNext;
_d_uartInBufferTop = _q_uartInBufferTop;
_d_uartInHold = _q_uartInHold;
_d_uartOutBuffer_wenable0 = _q_uartOutBuffer_wenable0;
_d_uartOutBuffer_addr0 = _q_uartOutBuffer_addr0;
_d_uartOutBuffer_wenable1 = _q_uartOutBuffer_wenable1;
_d_uartOutBuffer_wdata1 = _q_uartOutBuffer_wdata1;
_d_uartOutBuffer_addr1 = _q_uartOutBuffer_addr1;
_d_uartOutBufferNext = _q_uartOutBufferNext;
_d_uartOutBufferTop = _q_uartOutBufferTop;
_d_newuartOutBufferTop = _q_newuartOutBufferTop;
_d_uartOutHold = _q_uartOutHold;
_d_led = _q_led;
_d_uart_tx_data = _q_uart_tx_data;
_d_uart_tx_valid = _q_uart_tx_valid;
_d_sdram_cle = _q_sdram_cle;
_d_sdram_dqm = _q_sdram_dqm;
_d_sdram_cs = _q_sdram_cs;
_d_sdram_we = _q_sdram_we;
_d_sdram_cas = _q_sdram_cas;
_d_sdram_ras = _q_sdram_ras;
_d_sdram_ba = _q_sdram_ba;
_d_sdram_a = _q_sdram_a;
_d_sdram_clk = _q_sdram_clk;
_d_display_gpu_x = _q_display_gpu_x;
_d_display_gpu_y = _q_display_gpu_y;
_d_display_gpu_dotset = _q_display_gpu_dotset;
_d_display_gpu_write = _q_display_gpu_write;
_d_display_tpu_x = _q_display_tpu_x;
_d_display_tpu_y = _q_display_tpu_y;
_d_display_tpu_set = _q_display_tpu_set;
_d_display_tpu_write = _q_display_tpu_write;
_d_index = _q_index;
_vga_driver_run = 1;
_display_run = 1;
// _always_pre
_d_dstack_wenable = 0;
_d_rstack_wenable = 0;
_d_uartInBuffer_wenable0 = 0;
_d_uartInBuffer_wenable1 = 1;
_d_uartInBuffer_addr0 = _q_uartInBufferNext;
_d_uartInBuffer_addr1 = _q_uartInBufferTop;
_d_uartOutBuffer_wenable0 = 0;
_d_uartOutBuffer_wenable1 = 1;
_d_uartOutBuffer_addr0 = _q_uartOutBufferNext;
_d_uartOutBuffer_addr1 = _q_uartOutBufferTop;
_d_sdram_cle = 1'bz;
_d_sdram_dqm = 1'bz;
_d_sdram_cs = 1'bz;
_d_sdram_we = 1'bz;
_d_sdram_cas = 1'bz;
_d_sdram_ras = 1'bz;
_d_sdram_ba = 2'bz;
_d_sdram_a = 13'bz;
_d_sdram_clk = 1'bz;
_d_index = 7;
case (_q_index)
0: begin
// _top
// var inits
_d_pc = 0;
_d_dstack_wenable = 0;
_d_dstack_wdata = 0;
_d_dstack_addr = 0;
_d_stackTop = 0;
_d_dsp = 0;
_d_rstack_wenable = 0;
_d_rstack_wdata = 0;
_d_rstack_addr = 0;
_d_rsp = 0;
_d_rom_addr = 0;
_d_ram_wenable0 = 0;
_d_ram_wdata0 = 0;
_d_ram_addr0 = 0;
_d_ram_wenable1 = 0;
_d_ram_addr1 = 0;
_d_CYCLE = 0;
_d_INIT = 0;
_d_copyaddress = 0;
_d_bramREAD = 0;
_d_uartInBuffer_wenable0 = 0;
_d_uartInBuffer_addr0 = 0;
_d_uartInBuffer_wenable1 = 0;
_d_uartInBuffer_wdata1 = 0;
_d_uartInBuffer_addr1 = 0;
_d_uartInBufferNext = 0;
_d_uartInBufferTop = 0;
_d_uartInHold = 1;
_d_uartOutBuffer_wenable0 = 0;
_d_uartOutBuffer_addr0 = 0;
_d_uartOutBuffer_wenable1 = 0;
_d_uartOutBuffer_wdata1 = 0;
_d_uartOutBuffer_addr1 = 0;
_d_uartOutBufferNext = 0;
_d_uartOutBufferTop = 0;
_d_newuartOutBufferTop = 0;
_d_uartOutHold = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (_q_INIT==0) begin
// __block_2
// __block_4
  case (_q_CYCLE)
  0: begin
// __block_6_case
// __block_7
_d_ram_addr0 = _q_copyaddress;
_d_ram_wdata0 = 0;
_d_ram_wenable0 = 1;
// __block_8
  end
  1: begin
// __block_9_case
// __block_10
_d_copyaddress = _q_copyaddress+1;
_d_ram_wenable0 = 0;
// __block_11
  end
  4: begin
// __block_12_case
// __block_13
if (_q_copyaddress==32768) begin
// __block_14
// __block_16
_d_INIT = 1;
_d_copyaddress = 0;
// __block_17
end else begin
// __block_15
end
// __block_18
// __block_19
  end
  default: begin
// __block_20_case
// __block_21
// __block_22
  end
endcase
// __block_5
_d_CYCLE = (_q_CYCLE==4)?0:_q_CYCLE+1;
// __block_23
_d_index = 1;
end else begin
_d_index = 3;
end
end
3: begin
// __while__block_24
if (_q_INIT==1) begin
// __block_25
// __block_27
  case (_q_CYCLE)
  0: begin
// __block_29_case
// __block_30
_d_rom_addr = _q_copyaddress;
// __block_31
  end
  1: begin
// __block_32_case
// __block_33
_d_bramREAD = _w_mem_rom_rdata;
// __block_34
  end
  2: begin
// __block_35_case
// __block_36
_d_ram_addr0 = _q_copyaddress;
_d_ram_wdata0 = _q_bramREAD;
_d_ram_wenable0 = 1;
// __block_37
  end
  3: begin
// __block_38_case
// __block_39
_d_copyaddress = _q_copyaddress+1;
_d_ram_wenable0 = 0;
// __block_40
  end
  4: begin
// __block_41_case
// __block_42
if (_q_copyaddress==4096) begin
// __block_43
// __block_45
_d_INIT = 3;
_d_copyaddress = 0;
// __block_46
end else begin
// __block_44
end
// __block_47
// __block_48
  end
  default: begin
// __block_49_case
// __block_50
// __block_51
  end
endcase
// __block_28
_d_CYCLE = (_q_CYCLE==4)?0:_q_CYCLE+1;
// __block_52
_d_index = 3;
end else begin
_d_index = 5;
end
end
5: begin
// __while__block_53
if (_q_INIT==3) begin
// __block_54
// __block_56
  case (_q_uartInHold)
  0: begin
// __block_58_case
// __block_59
if (in_uart_rx_valid) begin
// __block_60
// __block_62
_d_uartInBuffer_wdata1 = in_uart_rx_data;
_d_uartInBufferTop = _q_uartInBufferTop+1;
_d_uartInHold = 1;
// __block_63
end else begin
// __block_61
end
// __block_64
// __block_65
  end
  1: begin
// __block_66_case
// __block_67
_d_uartInHold = (in_uart_rx_valid==0)?0:1;
// __block_68
  end
endcase
// __block_57
  case (_q_uartOutHold)
  0: begin
// __block_70_case
// __block_71
if (~(_q_uartOutBufferNext==_q_uartOutBufferTop)&~(in_uart_tx_busy)) begin
// __block_72
// __block_74
_d_uart_tx_data = _w_mem_uartOutBuffer_rdata0;
_d_uart_tx_valid = 1;
_d_uartOutHold = 1;
_d_uartOutBufferNext = _q_uartOutBufferNext+1;
// __block_75
end else begin
// __block_73
end
// __block_76
// __block_77
  end
  1: begin
// __block_78_case
// __block_79
if (~in_uart_tx_busy) begin
// __block_80
// __block_82
_d_uart_tx_valid = 0;
_d_uartOutHold = 0;
// __block_83
end else begin
// __block_81
end
// __block_84
// __block_85
  end
endcase
// __block_69
_d_uartOutBufferTop = _q_newuartOutBufferTop;
  case (_q_CYCLE)
  0: begin
// __block_87_case
// __block_88
_d_stackNext = _w_mem_dstack_rdata;
_d_rStackTop = _w_mem_rstack_rdata;
_d_ram_addr0 = _q_stackTop>>1;
_d_ram_wenable0 = 0;
_d_ram_addr1 = _q_pc;
_d_ram_wenable1 = 0;
// __block_89
  end
  1: begin
// __block_90_case
// __block_91
_d_memoryInput = _w_mem_ram_rdata0;
_d_instruction = _w_mem_ram_rdata1;
// __block_92
  end
  2: begin
// __block_93_case
// __block_94
if (_w_is_lit) begin
// __block_95
// __block_97
_d_newStackTop = _w_immediate;
_d_newPC = _w_pcPlusOne;
_d_newDSP = _q_dsp+1;
_d_newRSP = _q_rsp;
// __block_98
end else begin
// __block_96
// __block_99
  case (_q_instruction[13+:2])
  2'b00: begin
// __block_101_case
// __block_102
_d_newStackTop = _q_stackTop;
_d_newPC = _q_instruction[0+:13];
_d_newDSP = _q_dsp;
_d_newRSP = _q_rsp;
// __block_103
  end
  2'b01: begin
// __block_104_case
// __block_105
_d_newStackTop = _q_stackNext;
_d_newPC = (_q_stackTop==0)?_q_instruction[0+:13]:_w_pcPlusOne;
_d_newDSP = _q_dsp-1;
_d_newRSP = _q_rsp;
// __block_106
  end
  2'b10: begin
// __block_107_case
// __block_108
_d_newStackTop = _q_stackTop;
_d_newPC = _q_instruction[0+:13];
_d_newDSP = _q_dsp;
_d_newRSP = _q_rsp+1;
_d_rstackWData = _w_pcPlusOne<<1;
// __block_109
  end
  2'b11: begin
// __block_110_case
// __block_111
  case (_q_instruction[4+:1])
  1'b0: begin
// __block_113_case
// __block_114
  case (_q_instruction[8+:4])
  4'b0000: begin
// __block_116_case
// __block_117
_d_newStackTop = _q_stackTop;
// __block_118
  end
  4'b0001: begin
// __block_119_case
// __block_120
_d_newStackTop = _q_stackNext;
// __block_121
  end
  4'b0010: begin
// __block_122_case
// __block_123
_d_newStackTop = _q_stackTop+_q_stackNext;
// __block_124
  end
  4'b0011: begin
// __block_125_case
// __block_126
_d_newStackTop = _q_stackTop&_q_stackNext;
// __block_127
  end
  4'b0100: begin
// __block_128_case
// __block_129
_d_newStackTop = _q_stackTop|_q_stackNext;
// __block_130
  end
  4'b0101: begin
// __block_131_case
// __block_132
_d_newStackTop = _q_stackTop^_q_stackNext;
// __block_133
  end
  4'b0110: begin
// __block_134_case
// __block_135
_d_newStackTop = ~_q_stackTop;
// __block_136
  end
  4'b0111: begin
// __block_137_case
// __block_138
_d_newStackTop = {16{(_q_stackNext==_q_stackTop)}};
// __block_139
  end
  4'b1000: begin
// __block_140_case
// __block_141
_d_newStackTop = {16{($signed(_q_stackNext)<$signed(_q_stackTop))}};
// __block_142
  end
  4'b1001: begin
// __block_143_case
// __block_144
_d_newStackTop = _q_stackNext>>_q_stackTop[0+:4];
// __block_145
  end
  4'b1010: begin
// __block_146_case
// __block_147
_d_newStackTop = _q_stackTop-1;
// __block_148
  end
  4'b1011: begin
// __block_149_case
// __block_150
_d_newStackTop = _q_rStackTop;
// __block_151
  end
  4'b1100: begin
// __block_152_case
// __block_153
  case (_q_stackTop)
  16'hf000: begin
// __block_155_case
// __block_156
_d_newStackTop = {8'b0,_w_mem_uartInBuffer_rdata0};
_d_uartInBufferNext = _q_uartInBufferNext+1;
// __block_157
  end
  16'hf001: begin
// __block_158_case
// __block_159
_d_newStackTop = {14'b0,(_d_uartOutBufferTop+1==_d_uartOutBufferNext),~(_q_uartInBufferNext==_d_uartInBufferTop)};
// __block_160
  end
  16'hf002: begin
// __block_161_case
// __block_162
_d_newStackTop = _q_led;
// __block_163
  end
  16'hf003: begin
// __block_164_case
// __block_165
_d_newStackTop = {12'b0,in_buttons};
// __block_166
  end
  16'hf004: begin
// __block_167_case
// __block_168
_d_newStackTop = in_timer1hz;
// __block_169
  end
  default: begin
// __block_170_case
// __block_171
_d_newStackTop = _q_memoryInput;
// __block_172
  end
endcase
// __block_154
// __block_173
  end
  4'b1101: begin
// __block_174_case
// __block_175
_d_newStackTop = _q_stackNext<<_q_stackTop[0+:4];
// __block_176
  end
  4'b1110: begin
// __block_177_case
// __block_178
_d_newStackTop = {_q_rsp,_q_dsp};
// __block_179
  end
  4'b1111: begin
// __block_180_case
// __block_181
_d_newStackTop = {16{($unsigned(_q_stackNext)<$unsigned(_q_stackTop))}};
// __block_182
  end
endcase
// __block_115
// __block_183
  end
  1'b1: begin
// __block_184_case
// __block_185
  case (_q_instruction[8+:4])
  4'b0000: begin
// __block_187_case
// __block_188
_d_newStackTop = {16{(_q_stackTop==0)}};
// __block_189
  end
  4'b0001: begin
// __block_190_case
// __block_191
_d_newStackTop = ~{16{(_q_stackTop==0)}};
// __block_192
  end
  4'b0010: begin
// __block_193_case
// __block_194
_d_newStackTop = ~{16{(_q_stackNext==_q_stackTop)}};
// __block_195
  end
  4'b0011: begin
// __block_196_case
// __block_197
_d_newStackTop = _q_stackTop+1;
// __block_198
  end
  4'b0100: begin
// __block_199_case
// __block_200
_d_newStackTop = _q_stackTop<<1;
// __block_201
  end
  4'b0101: begin
// __block_202_case
// __block_203
_d_newStackTop = _q_stackTop>>1;
// __block_204
  end
  4'b0110: begin
// __block_205_case
// __block_206
_d_newStackTop = {16{($signed(_q_stackNext)>$signed(_q_stackTop))}};
// __block_207
  end
  4'b0111: begin
// __block_208_case
// __block_209
_d_newStackTop = {16{($unsigned(_q_stackNext)>$unsigned(_q_stackTop))}};
// __block_210
  end
  4'b1000: begin
// __block_211_case
// __block_212
_d_newStackTop = {16{($signed(_q_stackTop)<$signed(0))}};
// __block_213
  end
  4'b1001: begin
// __block_214_case
// __block_215
_d_newStackTop = {16{($signed(_q_stackTop)>$signed(0))}};
// __block_216
  end
  4'b1010: begin
// __block_217_case
// __block_218
_d_newStackTop = ($signed(_q_stackTop)<$signed(0))?-_q_stackTop:_q_stackTop;
// __block_219
  end
  4'b1011: begin
// __block_220_case
// __block_221
_d_newStackTop = ($signed(_q_stackNext)>$signed(_q_stackTop))?_q_stackNext:_q_stackTop;
// __block_222
  end
  4'b1100: begin
// __block_223_case
// __block_224
_d_newStackTop = ($signed(_q_stackNext)<$signed(_q_stackTop))?_q_stackNext:_q_stackTop;
// __block_225
  end
  4'b1101: begin
// __block_226_case
// __block_227
_d_newStackTop = -_q_stackTop;
// __block_228
  end
  4'b1110: begin
// __block_229_case
// __block_230
_d_newStackTop = _q_stackNext-_q_stackTop;
// __block_231
  end
  4'b1111: begin
// __block_232_case
// __block_233
_d_newStackTop = {16{($signed(_q_stackNext)>=$signed(_q_stackTop))}};
// __block_234
  end
endcase
// __block_186
// __block_235
  end
endcase
// __block_112
_d_newDSP = _q_dsp+_w_ddelta;
_d_newRSP = _q_rsp+_w_rdelta;
_d_rstackWData = _q_stackTop;
_d_newPC = (_q_instruction[12+:1])?_q_rStackTop>>1:_w_pcPlusOne;
if (_q_instruction[5+:1]) begin
// __block_236
// __block_238
  case (_q_stackTop)
  default: begin
// __block_240_case
// __block_241
_d_ram_addr0 = _q_stackTop>>1;
_d_ram_wdata0 = _q_stackNext;
_d_ram_wenable0 = 1;
// __block_242
  end
  16'hf000: begin
// __block_243_case
// __block_244
_d_uartOutBuffer_wdata1 = _q_stackNext[0+:8];
_d_newuartOutBufferTop = _d_uartOutBufferTop+1;
// __block_245
  end
  16'hf002: begin
// __block_246_case
// __block_247
_d_led = _q_stackNext;
// __block_248
  end
  16'hff00: begin
// __block_249_case
// __block_250
_d_display_gpu_x = _q_stackNext;
// __block_251
  end
  16'hff01: begin
// __block_252_case
// __block_253
_d_display_gpu_y = _q_stackNext;
// __block_254
  end
  16'hff02: begin
// __block_255_case
// __block_256
_d_display_gpu_dotset = _q_stackNext;
_d_display_gpu_write = 1;
// __block_257
  end
  16'hff10: begin
// __block_258_case
// __block_259
_d_display_tpu_x = _q_stackNext;
// __block_260
  end
  16'hff11: begin
// __block_261_case
// __block_262
_d_display_tpu_y = _q_stackNext;
// __block_263
  end
  16'hff12: begin
// __block_264_case
// __block_265
_d_display_tpu_set = _q_stackNext;
_d_display_tpu_write = 1;
// __block_266
  end
  16'hff13: begin
// __block_267_case
// __block_268
_d_display_tpu_set = _q_stackNext;
_d_display_tpu_write = 2;
// __block_269
  end
  16'hff14: begin
// __block_270_case
// __block_271
_d_display_tpu_set = _q_stackNext;
_d_display_tpu_write = 3;
// __block_272
  end
endcase
// __block_239
// __block_273
end else begin
// __block_237
end
// __block_274
// __block_275
  end
endcase
// __block_100
// __block_276
end
// __block_277
// __block_278
  end
  3: begin
// __block_279_case
// __block_280
if (_w_dstackWrite) begin
// __block_281
// __block_283
_d_dstack_wenable = 1;
_d_dstack_addr = _q_newDSP;
_d_dstack_wdata = _q_stackTop;
// __block_284
end else begin
// __block_282
end
// __block_285
if (_w_rstackWrite) begin
// __block_286
// __block_288
_d_rstack_wenable = 1;
_d_rstack_addr = _q_newRSP;
_d_rstack_wdata = _q_rstackWData;
// __block_289
end else begin
// __block_287
end
// __block_290
// __block_291
  end
  4: begin
// __block_292_case
// __block_293
_d_dsp = _q_newDSP;
_d_pc = _q_newPC;
_d_stackTop = _q_newStackTop;
_d_rsp = _q_newRSP;
_d_dstack_addr = _q_newDSP;
_d_rstack_addr = _q_newRSP;
_d_ram_wenable0 = 0;
_d_display_gpu_write = 0;
_d_display_tpu_write = 0;
// __block_294
  end
  default: begin
// __block_295_case
// __block_296
// __block_297
  end
endcase
// __block_86
_d_CYCLE = (_q_CYCLE==4)?0:_q_CYCLE+1;
// __block_298
_d_index = 5;
end else begin
_d_index = 6;
end
end
6: begin
// __block_55
_d_index = 7;
end
7: begin // end of main
end
default: begin 
_d_index = 7;
 end
endcase
end
endmodule

