`define HDMI 1
`define UART 1
`define BUTTONS 1
`define AUDIO 1
`define ULX3S 1
`default_nettype none

module top(
  // basic
  output [7:0] leds,
  // buttons
  input  [6:0] btns,
`ifdef SDRAM
  // sdram
  output sdram_clk,
  output sdram_cke,
  output [1:0]  sdram_dqm,
  output sdram_csn,
  output sdram_wen,
  output sdram_casn,
  output sdram_rasn,
  output [1:0]  sdram_ba,
  output [12:0] sdram_a,
  inout  [15:0] sdram_d,
`endif  
`ifdef AUDIO
  output [3:0] audio_l,
  output [3:0] audio_r,
`endif  
`ifdef OLED  
  // oled
  output  oled_clk,
  output  oled_mosi,
  output  oled_dc,
  output  oled_resn,
  output  oled_csn,
`endif  
`ifdef SDCARD
  // sdcard
  output  sd_clk,
  output  sd_csn,
  output  sd_mosi,
  input   sd_miso,
`endif  
`ifdef GPIO
  // gpio
  output [27:0] gp,
  input  [27:0] gn,
`endif  
`ifdef VGA
  // vga
  output [27:0] gp,
  input  [27:0] gn,
`endif  
`ifdef HDMI
  // hdmi
  output [3:0]  gpdi_dp, // {clock,R,G,B}
  output [3:0]  gpdi_dn,
`endif  
`ifdef UART
  // uart
  output  ftdi_rxd,
  input   ftdi_txd,
`endif
`ifdef UART2
  // uart2
`endif
  input  clk_25mhz
  );

wire [7:0]  __main_out_leds;

`ifdef OLED
wire        __main_oled_clk;
wire        __main_oled_mosi;
wire        __main_oled_dc;
wire        __main_oled_resn;
wire        __main_oled_csn;
`endif

`ifdef SDRAM
wire        __main_out_sdram_clk;
wire        __main_out_sdram_cle;
wire [1:0]  __main_out_sdram_dqm;
wire        __main_out_sdram_cs;
wire        __main_out_sdram_we;
wire        __main_out_sdram_cas;
wire        __main_out_sdram_ras;
wire [1:0]  __main_out_sdram_ba;
wire [12:0] __main_out_sdram_a;
`endif

`ifdef UART2
`ifndef GPIO
`error_UART2_needs_GPIO
`endif
`endif

`ifdef UART
wire        __main_out_uart_tx;
`endif

`ifdef VGA
wire        __main_out_vga_hs;
wire        __main_out_vga_vs;
wire [5:0]  __main_out_vga_r;
wire [5:0]  __main_out_vga_g;
wire [5:0]  __main_out_vga_b;
`endif

`ifdef SDCARD
wire        __main_sd_clk;
wire        __main_sd_csn;
wire        __main_sd_mosi;
`endif

`ifdef HDMI
wire [3:0]  __main_out_gpdi_dp;
wire [3:0]  __main_out_gpdi_dn;
`endif

`ifdef AUDIO
wire [3:0]  __main_out_audio_l;
wire [3:0]  __main_out_audio_r;
`endif

wire ready = btns[0];

reg [31:0] RST_d;
reg [31:0] RST_q;

always @* begin
  RST_d = RST_q >> 1;
end

always @(posedge clk_25mhz) begin
  if (ready) begin
    RST_q <= RST_d;
  end else begin
    RST_q <= 32'b111111111111111111111111111111;
  end
end

wire run_main;
assign run_main = 1'b1;

M_main __main(
  .reset         (RST_q[0]),
  .in_run        (run_main),
  .out_leds      (__main_out_leds),
`ifdef BUTTONS  
  .in_btns       (btns),
`endif
`ifdef SDRAM
  .inout_sdram_dq(sdram_d),
  .out_sdram_clk (__main_out_sdram_clk),
  .out_sdram_cle (__main_out_sdram_cle),
  .out_sdram_dqm (__main_out_sdram_dqm),
  .out_sdram_cs  (__main_out_sdram_cs),
  .out_sdram_we  (__main_out_sdram_we),
  .out_sdram_cas (__main_out_sdram_cas),
  .out_sdram_ras (__main_out_sdram_ras),
  .out_sdram_ba  (__main_out_sdram_ba),
  .out_sdram_a   (__main_out_sdram_a),
`endif  
`ifdef SDCARD
  .out_sd_csn    (__main_sd_csn),
  .out_sd_clk    (__main_sd_clk),
  .out_sd_mosi   (__main_sd_mosi),
  .in_sd_miso    (sd_miso),
`endif  
`ifdef AUDIO
  .out_audio_l  (__main_out_audio_l),
  .out_audio_r  (__main_out_audio_r),
`endif  
`ifdef OLED
  .out_oled_clk (__main_oled_clk),
  .out_oled_mosi(__main_oled_mosi),
  .out_oled_dc  (__main_oled_dc),
  .out_oled_resn(__main_oled_resn),
  .out_oled_csn (__main_oled_csn),
`endif 
`ifdef GPIO
`ifdef UART2
  .out_gp       (gp[27:1]),
  .in_gn        (gn[27:1]),
  .out_uart2_tx (gp[0]),
  .in_uart2_rx  (gn[0]),
`else
  .out_gp       (gp),
  .in_gn        (gn),
`endif  
`endif  
`ifdef UART
  .out_uart_tx  (__main_out_uart_tx),
  .in_uart_rx   (ftdi_txd),
`endif  
`ifdef VGA
  .out_video_hs (__main_out_vga_hs),
  .out_video_vs (__main_out_vga_vs),
  .out_video_r  (__main_out_vga_r),
  .out_video_g  (__main_out_vga_g),
  .out_video_b  (__main_out_vga_b),  
`endif  
`ifdef HDMI
  .out_gpdi_dp  (__main_out_gpdi_dp),
  .out_gpdi_dn  (__main_out_gpdi_dn),
`endif
  .clock         (clk_25mhz)
);

assign leds          = __main_out_leds;

`ifdef SDRAM
assign sdram_clk     = __main_out_sdram_clk;
assign sdram_cke     = __main_out_sdram_cle;
assign sdram_dqm     = __main_out_sdram_dqm;
assign sdram_csn     = __main_out_sdram_cs;
assign sdram_wen     = __main_out_sdram_we;
assign sdram_casn    = __main_out_sdram_cas;
assign sdram_rasn    = __main_out_sdram_ras;
assign sdram_ba      = __main_out_sdram_ba;
assign sdram_a       = __main_out_sdram_a;
`endif

`ifdef AUDIO
assign audio_l       = __main_out_audio_l;
assign audio_r       = __main_out_audio_r;
`endif  

`ifdef VGA
assign gp[0]         = __main_out_vga_vs;
assign gp[1]         = __main_out_vga_hs;
assign gp[2]         = __main_out_vga_r[5];
assign gp[3]         = __main_out_vga_r[4];
assign gp[4]         = __main_out_vga_r[3];
assign gp[5]         = __main_out_vga_r[2];
assign gp[6]         = __main_out_vga_r[1];
assign gp[7]         = __main_out_vga_r[0];
assign gp[8]         = __main_out_vga_g[5];
assign gp[9]         = __main_out_vga_g[4];
assign gp[10]        = __main_out_vga_g[3];
assign gp[11]        = __main_out_vga_g[2];
assign gp[12]        = __main_out_vga_g[1];
assign gp[13]        = __main_out_vga_g[0];
assign gp[14]        = __main_out_vga_b[0];
assign gp[15]        = __main_out_vga_b[1];
assign gp[16]        = __main_out_vga_b[2];
assign gp[17]        = __main_out_vga_b[3];
assign gp[18]        = __main_out_vga_b[4];
assign gp[19]        = __main_out_vga_b[5];
`endif

`ifdef SDCARD
assign sd_clk        = __main_sd_clk;
assign sd_csn        = __main_sd_csn;
assign sd_mosi       = __main_sd_mosi;
`endif

`ifdef OLED
assign oled_clk      = __main_oled_clk;
assign oled_mosi     = __main_oled_mosi;
assign oled_dc       = __main_oled_dc;
assign oled_resn     = __main_oled_resn;
assign oled_csn      = __main_oled_csn;
`endif

`ifdef UART
assign ftdi_rxd      = __main_out_uart_tx;
`endif  

`ifdef HDMI
assign gpdi_dp       = __main_out_gpdi_dp;
assign gpdi_dn       = __main_out_gpdi_dn;
`endif

endmodule

module hdmi_clock (
        input  clk,           //  25 MHz
        output half_hdmi_clk  // 125 MHz
    );

`ifdef MOJO

`else

`ifdef DE10NANO

`else

`ifdef ULX3S

wire clkfb;
wire clkos;
wire clkout0;
wire clkout2;
wire locked;

(* ICP_CURRENT="12" *) (* LPF_RESISTOR="8" *) (* MFG_ENABLE_FILTEROPAMP="1" *) (* MFG_GMCREF_SEL="2" *)
EHXPLLL #(
        .PLLRST_ENA("DISABLED"),
        .INTFB_WAKE("DISABLED"),
        .STDBY_ENABLE("DISABLED"),
        .DPHASE_SOURCE("DISABLED"),
        .CLKOP_FPHASE(0),
        .CLKOP_CPHASE(0),
        .OUTDIVIDER_MUXA("DIVA"),
        .CLKOP_ENABLE("ENABLED"),
        .CLKOP_DIV(2),
        .CLKOS_ENABLE("ENABLED"),
        .CLKOS_DIV(4),
        .CLKOS_CPHASE(0),
        .CLKOS_FPHASE(0),
        .CLKOS2_ENABLE("ENABLED"),
        .CLKOS2_DIV(20),
        .CLKOS2_CPHASE(0),
        .CLKOS2_FPHASE(0),
        .CLKFB_DIV(10),
        .CLKI_DIV(1),
        .FEEDBK_PATH("INT_OP")
    ) pll_i (
        .CLKI(clk),
        .CLKFB(clkfb),
        .CLKINTFB(clkfb),
        .CLKOP(clkout0), // 250
        .CLKOS(half_hdmi_clk),  // 125
        .CLKOS2(clkout2), // 25
        .RST(1'b0),
        .STDBY(1'b0),
        .PHASESEL0(1'b0),
        .PHASESEL1(1'b0),
        .PHASEDIR(1'b0),
        .PHASESTEP(1'b0),
        .PLLWAKESYNC(1'b0),
        .ENCLKOP(1'b0),
        .LOCK(locked)
	);

`else

`ifdef ICARUS

reg genclk;

initial begin
  genclk = 1'b0;
  forever #4 genclk = ~genclk;   // generates a 125 MHz clock
end

assign half_hdmi_clk = genclk;

`endif
    
`endif
`endif
`endif
    
endmodule


// @sylefeb differential pair for HDMI, outputting dual rate
//
// see also https://github.com/lawrie/ulx3s_examples/blob/master/hdmi/fake_differential.v

module differential_pair(
        input   clock,
        input   [1:0] pos,
        input   [1:0] neg,
        output  out_pin_pos,
        output  out_pin_neg
    );

`ifdef ULX3S

ODDRX1F ddr_pos
      (
        .D0(pos[0]),
        .D1(pos[1]),
        .Q(out_pin_pos),
        .SCLK(clock),
        .RST(0)
      );

ODDRX1F ddr_neg
      (
        .D0(neg[0]),
        .D1(neg[1]),
        .Q(out_pin_neg),
        .SCLK(clock),
        .RST(0)
      );

`else

`ifdef ICARUS

assign out_pin_pos = pos[0];
assign out_pin_neg = neg[0];

`endif

`endif

endmodule


module hdmi_differential_pairs(
        input   clock,
        input   [7:0] pos,
        input   [7:0] neg,
        output  [3:0] out_pos,
        output  [3:0] out_neg
    );

  differential_pair rp(
    .clock(clock),
    .pos(pos[0+:2]),
    .neg(neg[0+:2]),
    .out_pin_pos(out_pos[2+:1]),
    .out_pin_neg(out_neg[2+:1])
  );

  differential_pair gp(
    .clock(clock),
    .pos(pos[2+:2]),
    .neg(neg[2+:2]),
    .out_pin_pos(out_pos[1+:1]),
    .out_pin_neg(out_neg[1+:1])
  );

  differential_pair bp(
    .clock(clock),
    .pos(pos[4+:2]),
    .neg(neg[4+:2]),
    .out_pin_pos(out_pos[0+:1]),
    .out_pin_neg(out_neg[0+:1])
  );

  differential_pair cp(
    .clock(clock),
    .pos(pos[6+:2]),
    .neg(neg[6+:2]),
    .out_pin_pos(out_pos[3+:1]),
    .out_pin_neg(out_neg[3+:1])
  );

endmodule


// diamond 3.7 accepts this PLL
// diamond 3.8-3.9 is untested
// diamond 3.10 or higher is likely to abort with error about unable to use feedback signal
// cause of this could be from wrong CPHASE/FPHASE parameters
module ulx3s_clk_50_25
(
    input clkin, // 25 MHz, 0 deg
    output clkout0, // 50 MHz, 0 deg
    output clkout1, // 25 MHz, 0 deg
    output locked
);
(* FREQUENCY_PIN_CLKI="25" *)
(* FREQUENCY_PIN_CLKOP="50" *)
(* FREQUENCY_PIN_CLKOS="25" *)
(* ICP_CURRENT="12" *) (* LPF_RESISTOR="8" *) (* MFG_ENABLE_FILTEROPAMP="1" *) (* MFG_GMCREF_SEL="2" *)
EHXPLLL #(
        .PLLRST_ENA("DISABLED"),
        .INTFB_WAKE("DISABLED"),
        .STDBY_ENABLE("DISABLED"),
        .DPHASE_SOURCE("DISABLED"),
        .OUTDIVIDER_MUXA("DIVA"),
        .OUTDIVIDER_MUXB("DIVB"),
        .OUTDIVIDER_MUXC("DIVC"),
        .OUTDIVIDER_MUXD("DIVD"),
        .CLKI_DIV(1),
        .CLKOP_ENABLE("ENABLED"),
        .CLKOP_DIV(12),
        .CLKOP_CPHASE(5),
        .CLKOP_FPHASE(0),
        .CLKOS_ENABLE("ENABLED"),
        .CLKOS_DIV(24),
        .CLKOS_CPHASE(5),
        .CLKOS_FPHASE(0),
        .FEEDBK_PATH("CLKOP"),
        .CLKFB_DIV(2)
    ) pll_i (
        .RST(1'b0),
        .STDBY(1'b0),
        .CLKI(clkin),
        .CLKOP(clkout0),
        .CLKOS(clkout1),
        .CLKFB(clkout0),
        .CLKINTFB(),
        .PHASESEL0(1'b0),
        .PHASESEL1(1'b0),
        .PHASEDIR(1'b1),
        .PHASESTEP(1'b1),
        .PHASELOADREG(1'b1),
        .PLLWAKESYNC(1'b0),
        .ENCLKOP(1'b0),
        .LOCK(locked)
	);
endmodule


module reset_conditioner (
    input rcclk,
    input in,
    output reg out
  );  
  reg [7:0] counter_d,counter_q;
  always @* begin
    counter_d = counter_q;
    if (counter_q == 0) begin
      out = 0;
    end else begin
      out = 1;
      counter_d = counter_q + 1;
    end
  end  
  always @(posedge rcclk) begin
    if (in == 1'b1) begin
      counter_q <= 1;
    end else begin
      counter_q <= counter_d;
    end
  end 
endmodule 


module M_tmds_encoder (
in_data,
in_ctrl,
in_data_or_ctrl,
out_tmds,
reset,
out_clock,
clock
);
input  [7:0] in_data;
input  [1:0] in_ctrl;
input  [0:0] in_data_or_ctrl;
output  [9:0] out_tmds;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [3:0] _w_num_ones;
wire signed [4:0] _w_diff_ones_zeros;
wire signed [0:0] _w_xored1;
wire signed [0:0] _w_xored2;
wire signed [0:0] _w_xored3;
wire signed [0:0] _w_xored4;
wire signed [0:0] _w_xored5;
wire signed [0:0] _w_xored6;
wire signed [0:0] _w_xored7;
wire signed [0:0] _w_xnored1;
wire signed [0:0] _w_xnored2;
wire signed [0:0] _w_xnored3;
wire signed [0:0] _w_xnored4;
wire signed [0:0] _w_xnored5;
wire signed [0:0] _w_xnored6;
wire signed [0:0] _w_xnored7;

reg  [8:0] _d_q_m;
reg  [8:0] _q_q_m;
reg signed [4:0] _d_dc_bias;
reg signed [4:0] _q_dc_bias;
reg  [9:0] _d_tmds,_q_tmds;
assign out_tmds = _q_tmds;

always @(posedge clock) begin
  if (reset) begin
_q_q_m <= 0;
_q_dc_bias <= 0;
  end else begin
_q_q_m <= _d_q_m;
_q_dc_bias <= _d_dc_bias;
_q_tmds <= _d_tmds;
  end
end



assign _w_xnored7 = ~(in_data[7+:1]^_w_xnored6);
assign _w_xnored5 = ~(in_data[5+:1]^_w_xnored4);
assign _w_xnored1 = ~(in_data[1+:1]^in_data[0+:1]);
assign _w_xored1 = in_data[1+:1]^in_data[0+:1];
assign _w_xored2 = in_data[2+:1]^_w_xored1;
assign _w_xored3 = in_data[3+:1]^_w_xored2;
assign _w_xored4 = in_data[4+:1]^_w_xored3;
assign _w_xnored6 = ~(in_data[6+:1]^_w_xnored5);
assign _w_xored5 = in_data[5+:1]^_w_xored4;
assign _w_xored6 = in_data[6+:1]^_w_xored5;
assign _w_xored7 = in_data[7+:1]^_w_xored6;
assign _w_xnored2 = ~(in_data[2+:1]^_w_xnored1);
assign _w_diff_ones_zeros = _d_q_m[0+:1]+_d_q_m[1+:1]+_d_q_m[2+:1]+_d_q_m[3+:1]+_d_q_m[4+:1]+_d_q_m[5+:1]+_d_q_m[6+:1]+_d_q_m[7+:1]-6'd4;
assign _w_xnored3 = ~(in_data[3+:1]^_w_xnored2);
assign _w_num_ones = in_data[0+:1]+in_data[1+:1]+in_data[2+:1]+in_data[3+:1]+in_data[4+:1]+in_data[5+:1]+in_data[6+:1]+in_data[7+:1];
assign _w_xnored4 = ~(in_data[4+:1]^_w_xnored3);

always @* begin
_d_q_m = _q_q_m;
_d_dc_bias = _q_dc_bias;
_d_tmds = _q_tmds;
// _always_pre
if ((_w_num_ones>4)||(_w_num_ones==4&&in_data[0+:1]==0)) begin
// __block_1
// __block_3
_d_q_m = {1'b0,{_w_xnored7,_w_xnored6,_w_xnored5,_w_xnored4,_w_xnored3,_w_xnored2,_w_xnored1},in_data[0+:1]};
// __block_4
end else begin
// __block_2
// __block_5
_d_q_m = {1'b1,{_w_xored7,_w_xored6,_w_xored5,_w_xored4,_w_xored3,_w_xored2,_w_xored1},in_data[0+:1]};
// __block_6
end
// __block_7
if (in_data_or_ctrl) begin
// __block_8
// __block_10
if (_q_dc_bias==0||_w_diff_ones_zeros==0) begin
// __block_11
// __block_13
_d_tmds = {~_d_q_m[8+:1],_d_q_m[8+:1],(_d_q_m[8+:1]?_d_q_m[0+:8]:~_d_q_m[0+:8])};
if (_d_q_m[8+:1]==0) begin
// __block_14
// __block_16
_d_dc_bias = _q_dc_bias-_w_diff_ones_zeros;
// __block_17
end else begin
// __block_15
// __block_18
_d_dc_bias = _q_dc_bias+_w_diff_ones_zeros;
// __block_19
end
// __block_20
// __block_21
end else begin
// __block_12
// __block_22
if ((_q_dc_bias>0&&_w_diff_ones_zeros>0)||(_q_dc_bias<0&&_w_diff_ones_zeros<0)) begin
// __block_23
// __block_25
_d_tmds = {1'b1,_d_q_m[8+:1],~_d_q_m[0+:8]};
_d_dc_bias = _q_dc_bias+_d_q_m[8+:1]-_w_diff_ones_zeros;
// __block_26
end else begin
// __block_24
// __block_27
_d_tmds = {1'b0,_d_q_m};
_d_dc_bias = _q_dc_bias-(~_d_q_m[8+:1])+_w_diff_ones_zeros;
// __block_28
end
// __block_29
// __block_30
end
// __block_31
// __block_32
end else begin
// __block_9
// __block_33
  case (in_ctrl)
  2'b00: begin
// __block_35_case
// __block_36
_d_tmds = 10'b1101010100;
// __block_37
  end
  2'b01: begin
// __block_38_case
// __block_39
_d_tmds = 10'b0010101011;
// __block_40
  end
  2'b10: begin
// __block_41_case
// __block_42
_d_tmds = 10'b0101010100;
// __block_43
  end
  2'b11: begin
// __block_44_case
// __block_45
_d_tmds = 10'b1010101011;
// __block_46
  end
endcase
// __block_34
_d_dc_bias = 0;
// __block_47
end
// __block_48
end
endmodule


module M_hdmi_ddr_shifter (
in_data_r,
in_data_g,
in_data_b,
out_outbits,
reset,
out_clock,
clock
);
input  [9:0] in_data_r;
input  [9:0] in_data_g;
input  [9:0] in_data_b;
output  [7:0] out_outbits;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
reg  [1:0] _t_clkbits;

reg  [2:0] _d_mod5;
reg  [2:0] _q_mod5;
reg  [9:0] _d_shift_r;
reg  [9:0] _q_shift_r;
reg  [9:0] _d_shift_g;
reg  [9:0] _q_shift_g;
reg  [9:0] _d_shift_b;
reg  [9:0] _q_shift_b;
reg  [7:0] _d_outbits,_q_outbits;
assign out_outbits = _q_outbits;

always @(posedge clock) begin
  if (reset) begin
_q_mod5 <= 0;
_q_shift_r <= 0;
_q_shift_g <= 0;
_q_shift_b <= 0;
  end else begin
_q_mod5 <= _d_mod5;
_q_shift_r <= _d_shift_r;
_q_shift_g <= _d_shift_g;
_q_shift_b <= _d_shift_b;
_q_outbits <= _d_outbits;
  end
end




always @* begin
_d_mod5 = _q_mod5;
_d_shift_r = _q_shift_r;
_d_shift_g = _q_shift_g;
_d_shift_b = _q_shift_b;
_d_outbits = _q_outbits;
_t_clkbits = 0;
// _always_pre
_d_shift_r = (_q_mod5==0)?in_data_r:_q_shift_r[2+:8];
_d_shift_g = (_q_mod5==0)?in_data_g:_q_shift_g[2+:8];
_d_shift_b = (_q_mod5==0)?in_data_b:_q_shift_b[2+:8];
_t_clkbits = (_q_mod5[0+:2]<2)?2'b11:((_q_mod5>2)?2'b00:2'b01);
_d_outbits = {_t_clkbits,_d_shift_b[0+:2],_d_shift_g[0+:2],_d_shift_r[0+:2]};
_d_mod5 = (_q_mod5==4)?0:(_q_mod5+1);
end
endmodule


module M_hdmi (
in_red,
in_green,
in_blue,
out_x,
out_y,
out_active,
out_vblank,
out_gpdi_dp,
out_gpdi_dn,
reset,
out_clock,
clock
);
input  [7:0] in_red;
input  [7:0] in_green;
input  [7:0] in_blue;
output  [9:0] out_x;
output  [9:0] out_y;
output  [0:0] out_active;
output  [0:0] out_vblank;
output  [3:0] out_gpdi_dp;
output  [3:0] out_gpdi_dn;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire[3:0] _w_hdmi_out_out_pos;
wire[3:0] _w_hdmi_out_out_neg;
wire _w_pll_half_hdmi_clk;
wire  [9:0] _w_tmdsR_tmds;
wire  [9:0] _w_tmdsG_tmds;
wire  [9:0] _w_tmdsB_tmds;
wire  [7:0] _w_shift_outbits;
wire  [1:0] _c_null_ctrl;
assign _c_null_ctrl = 0;
reg  [0:0] _t_hsync;
reg  [0:0] _t_vsync;
wire  [7:0] _w_crgb_neg;

reg  [9:0] _d_cntx;
reg  [9:0] _q_cntx;
reg  [9:0] _d_cnty;
reg  [9:0] _q_cnty;
reg  [1:0] _d_sync_ctrl;
reg  [1:0] _q_sync_ctrl;
reg  [7:0] _d_latch_red;
reg  [7:0] _q_latch_red;
reg  [7:0] _d_latch_green;
reg  [7:0] _q_latch_green;
reg  [7:0] _d_latch_blue;
reg  [7:0] _q_latch_blue;
reg  [1:0] _d_prev_sync_ctrl;
reg  [1:0] _q_prev_sync_ctrl;
reg  [0:0] _d_prev_active;
reg  [0:0] _q_prev_active;
reg  [9:0] _d_x,_q_x;
reg  [9:0] _d_y,_q_y;
reg  [0:0] _d_active,_q_active;
reg  [0:0] _d_vblank,_q_vblank;
assign out_x = _q_x;
assign out_y = _q_y;
assign out_active = _q_active;
assign out_vblank = _q_vblank;
assign out_gpdi_dp = _w_hdmi_out_out_pos;
assign out_gpdi_dn = _w_hdmi_out_out_neg;

always @(posedge clock) begin
  if (reset) begin
_q_cntx <= 0;
_q_cnty <= 0;
_q_sync_ctrl <= 0;
_q_latch_red <= 0;
_q_latch_green <= 0;
_q_latch_blue <= 0;
_q_prev_sync_ctrl <= 0;
_q_prev_active <= 0;
  end else begin
_q_cntx <= _d_cntx;
_q_cnty <= _d_cnty;
_q_sync_ctrl <= _d_sync_ctrl;
_q_latch_red <= _d_latch_red;
_q_latch_green <= _d_latch_green;
_q_latch_blue <= _d_latch_blue;
_q_prev_sync_ctrl <= _d_prev_sync_ctrl;
_q_prev_active <= _d_prev_active;
_q_x <= _d_x;
_q_y <= _d_y;
_q_active <= _d_active;
_q_vblank <= _d_vblank;
  end
end


hdmi_differential_pairs _hdmi_out (
.clock(_w_pll_half_hdmi_clk),
.pos(_w_shift_outbits),
.neg(_w_crgb_neg),
.out_pos(_w_hdmi_out_out_pos),
.out_neg(_w_hdmi_out_out_neg)
);

hdmi_clock _pll (
.clk(clock),
.half_hdmi_clk(_w_pll_half_hdmi_clk)
);
M_tmds_encoder tmdsR (
.in_data(_q_latch_red),
.in_ctrl(_c_null_ctrl),
.in_data_or_ctrl(_q_prev_active),
.out_tmds(_w_tmdsR_tmds),
.reset(reset),
.clock(clock)
);
M_tmds_encoder tmdsG (
.in_data(_q_latch_green),
.in_ctrl(_c_null_ctrl),
.in_data_or_ctrl(_q_prev_active),
.out_tmds(_w_tmdsG_tmds),
.reset(reset),
.clock(clock)
);
M_tmds_encoder tmdsB (
.in_data(_q_latch_blue),
.in_ctrl(_q_prev_sync_ctrl),
.in_data_or_ctrl(_q_prev_active),
.out_tmds(_w_tmdsB_tmds),
.reset(reset),
.clock(clock)
);
M_hdmi_ddr_shifter shift (
.in_data_r(_w_tmdsR_tmds),
.in_data_g(_w_tmdsG_tmds),
.in_data_b(_w_tmdsB_tmds),
.out_outbits(_w_shift_outbits),
.reset(reset),
.clock(_w_pll_half_hdmi_clk)
);


assign _w_crgb_neg = ~_w_shift_outbits;

always @* begin
_d_cntx = _q_cntx;
_d_cnty = _q_cnty;
_d_sync_ctrl = _q_sync_ctrl;
_d_latch_red = _q_latch_red;
_d_latch_green = _q_latch_green;
_d_latch_blue = _q_latch_blue;
_d_prev_sync_ctrl = _q_prev_sync_ctrl;
_d_prev_active = _q_prev_active;
_d_x = _q_x;
_d_y = _q_y;
_d_active = _q_active;
_d_vblank = _q_vblank;
_t_hsync = 0;
_t_vsync = 0;
// _always_pre
_d_prev_sync_ctrl = _q_sync_ctrl;
_d_prev_active = _q_active;
_t_hsync = (_q_cntx>655)&&(_q_cntx<752);
_t_vsync = (_q_cnty>489)&&(_q_cnty<492);
_d_sync_ctrl = {_t_vsync,_t_hsync};
_d_active = (_q_cntx<640)&&(_q_cnty<480);
_d_vblank = (_q_cnty>=480);
_d_x = (_q_cntx<640)?_q_cntx:0;
_d_y = (_q_cnty>=480)?0:_q_cnty;
_d_cnty = (_q_cntx==799)?(_q_cnty==524?0:(_q_cnty+1)):_q_cnty;
_d_cntx = (_q_cntx==799)?0:(_q_cntx+1);
_d_latch_red = in_red;
_d_latch_green = in_green;
_d_latch_blue = in_blue;
end
endmodule


module M_uart_sender #(
parameter IO_DATA_IN_WIDTH=1,parameter IO_DATA_IN_SIGNED=0,parameter IO_DATA_IN_INIT=0,
parameter IO_DATA_IN_READY_WIDTH=1,parameter IO_DATA_IN_READY_SIGNED=0,parameter IO_DATA_IN_READY_INIT=0,
parameter IO_BUSY_WIDTH=1,parameter IO_BUSY_SIGNED=0,parameter IO_BUSY_INIT=0
) (
in_io_data_in,
in_io_data_in_ready,
out_io_busy,
out_uart_tx,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [IO_DATA_IN_WIDTH-1:0] in_io_data_in;
input  [IO_DATA_IN_READY_WIDTH-1:0] in_io_data_in_ready;
output  [IO_BUSY_WIDTH-1:0] out_io_busy;
output  [0:0] out_uart_tx;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [9:0] _c_interval;
assign _c_interval = 434;

reg  [9:0] _d_counter;
reg  [9:0] _q_counter;
reg  [10:0] _d_transmit;
reg  [10:0] _q_transmit;
reg  [IO_BUSY_WIDTH-1:0] _d_io_busy,_q_io_busy;
reg  [0:0] _d_uart_tx,_q_uart_tx;
reg  [0:0] _d_index,_q_index;
assign out_io_busy = _q_io_busy;
assign out_uart_tx = _q_uart_tx;
assign out_done = (_q_index == 1);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_counter <= 0;
_q_transmit <= 0;
_q_io_busy <= IO_BUSY_INIT;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_counter <= _d_counter;
_q_transmit <= _d_transmit;
_q_io_busy <= _d_io_busy;
_q_uart_tx <= _d_uart_tx;
_q_index <= _d_index;
  end
end




always @* begin
_d_counter = _q_counter;
_d_transmit = _q_transmit;
_d_io_busy = _q_io_busy;
_d_uart_tx = _q_uart_tx;
_d_index = _q_index;
// _always_pre
if (_q_transmit>1) begin
// __block_1
// __block_3
if (_q_counter==0) begin
// __block_4
// __block_6
_d_uart_tx = _q_transmit[0+:1];
_d_transmit = {1'b0,_q_transmit[1+:10]};
// __block_7
end else begin
// __block_5
end
// __block_8
_d_counter = (_q_counter==_c_interval)?0:(_q_counter+1);
// __block_9
end else begin
// __block_2
// __block_10
_d_uart_tx = 1;
_d_io_busy = 0;
if (in_io_data_in_ready) begin
// __block_11
// __block_13
_d_io_busy = 1;
_d_transmit = {1'b1,1'b0,in_io_data_in,1'b0};
// __block_14
end else begin
// __block_12
end
// __block_15
// __block_16
end
// __block_17
_d_index = 1;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_counter = 0;
_d_transmit = 0;
// --
_d_uart_tx = 1;
_d_index = 1;
end
1: begin // end of uart_sender
end
default: begin 
_d_index = 1;
 end
endcase
end
endmodule


module M_uart_receiver #(
parameter IO_DATA_OUT_WIDTH=1,parameter IO_DATA_OUT_SIGNED=0,parameter IO_DATA_OUT_INIT=0,
parameter IO_DATA_OUT_READY_WIDTH=1,parameter IO_DATA_OUT_READY_SIGNED=0,parameter IO_DATA_OUT_READY_INIT=0
) (
in_uart_rx,
out_io_data_out,
out_io_data_out_ready,
reset,
out_clock,
clock
);
input  [0:0] in_uart_rx;
output  [IO_DATA_OUT_WIDTH-1:0] out_io_data_out;
output  [IO_DATA_OUT_READY_WIDTH-1:0] out_io_data_out_ready;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [9:0] _c_interval;
assign _c_interval = 434;
wire  [9:0] _c_half_interval;
assign _c_half_interval = 217;

reg  [9:0] _d_counter;
reg  [9:0] _q_counter;
reg  [3:0] _d_receiving;
reg  [3:0] _q_receiving;
reg  [9:0] _d_received;
reg  [9:0] _q_received;
reg  [0:0] _d_latched_rx;
reg  [0:0] _q_latched_rx;
reg  [IO_DATA_OUT_WIDTH-1:0] _d_io_data_out,_q_io_data_out;
reg  [IO_DATA_OUT_READY_WIDTH-1:0] _d_io_data_out_ready,_q_io_data_out_ready;
assign out_io_data_out = _q_io_data_out;
assign out_io_data_out_ready = _q_io_data_out_ready;

always @(posedge clock) begin
  if (reset) begin
_q_counter <= 0;
_q_receiving <= 0;
_q_received <= 0;
_q_latched_rx <= 0;
_q_io_data_out <= IO_DATA_OUT_INIT;
_q_io_data_out_ready <= IO_DATA_OUT_READY_INIT;
  end else begin
_q_counter <= _d_counter;
_q_receiving <= _d_receiving;
_q_received <= _d_received;
_q_latched_rx <= _d_latched_rx;
_q_io_data_out <= _d_io_data_out;
_q_io_data_out_ready <= _d_io_data_out_ready;
  end
end




always @* begin
_d_counter = _q_counter;
_d_receiving = _q_receiving;
_d_received = _q_received;
_d_latched_rx = _q_latched_rx;
_d_io_data_out = _q_io_data_out;
_d_io_data_out_ready = _q_io_data_out_ready;
// _always_pre
_d_io_data_out_ready = 0;
if (_q_receiving==0) begin
// __block_1
// __block_3
if (_q_latched_rx==0) begin
// __block_4
// __block_6
_d_receiving = 10;
_d_received = 0;
_d_counter = _c_half_interval;
// __block_7
end else begin
// __block_5
end
// __block_8
// __block_9
end else begin
// __block_2
// __block_10
if (_q_counter==0) begin
// __block_11
// __block_13
_d_received = {_q_latched_rx,_q_received[1+:9]};
_d_receiving = _q_receiving-1;
_d_counter = _c_interval;
if (_d_receiving==0) begin
// __block_14
// __block_16
_d_io_data_out = _d_received[1+:8];
_d_io_data_out_ready = 1;
// __block_17
end else begin
// __block_15
end
// __block_18
// __block_19
end else begin
// __block_12
// __block_20
_d_counter = _q_counter-1;
// __block_21
end
// __block_22
// __block_23
end
// __block_24
_d_latched_rx = in_uart_rx;
end
endmodule


module M_multiplex_display (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_background_r,
in_background_g,
in_background_b,
in_tilemap_r,
in_tilemap_g,
in_tilemap_b,
in_tilemap_display,
in_lower_sprites_r,
in_lower_sprites_g,
in_lower_sprites_b,
in_lower_sprites_display,
in_bitmap_r,
in_bitmap_g,
in_bitmap_b,
in_bitmap_display,
in_upper_sprites_r,
in_upper_sprites_g,
in_upper_sprites_b,
in_upper_sprites_display,
in_character_map_r,
in_character_map_g,
in_character_map_b,
in_character_map_display,
in_terminal_r,
in_terminal_g,
in_terminal_b,
in_terminal_display,
out_pix_red,
out_pix_green,
out_pix_blue,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [1:0] in_background_r;
input  [1:0] in_background_g;
input  [1:0] in_background_b;
input  [1:0] in_tilemap_r;
input  [1:0] in_tilemap_g;
input  [1:0] in_tilemap_b;
input  [0:0] in_tilemap_display;
input  [1:0] in_lower_sprites_r;
input  [1:0] in_lower_sprites_g;
input  [1:0] in_lower_sprites_b;
input  [0:0] in_lower_sprites_display;
input  [1:0] in_bitmap_r;
input  [1:0] in_bitmap_g;
input  [1:0] in_bitmap_b;
input  [0:0] in_bitmap_display;
input  [1:0] in_upper_sprites_r;
input  [1:0] in_upper_sprites_g;
input  [1:0] in_upper_sprites_b;
input  [0:0] in_upper_sprites_display;
input  [1:0] in_character_map_r;
input  [1:0] in_character_map_g;
input  [1:0] in_character_map_b;
input  [0:0] in_character_map_display;
input  [1:0] in_terminal_r;
input  [1:0] in_terminal_g;
input  [1:0] in_terminal_b;
input  [0:0] in_terminal_display;
output  [7:0] out_pix_red;
output  [7:0] out_pix_green;
output  [7:0] out_pix_blue;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [7:0] _w_RED_pix;
wire _w_RED_done;
wire  [7:0] _w_GREEN_pix;
wire _w_GREEN_done;
wire  [7:0] _w_BLUE_pix;
wire _w_BLUE_done;

reg  [7:0] _d_pix_red,_q_pix_red;
reg  [7:0] _d_pix_green,_q_pix_green;
reg  [7:0] _d_pix_blue,_q_pix_blue;
reg  [1:0] _d_index,_q_index;
reg  _RED_run;
reg  _GREEN_run;
reg  _BLUE_run;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_index <= _d_index;
  end
end

M_expandcolour RED (
.in_terminal_display(in_terminal_display),
.in_terminal(in_terminal_r),
.in_character_map_display(in_character_map_display),
.in_character_map(in_character_map_r),
.in_upper_sprites_display(in_upper_sprites_display),
.in_upper_sprites(in_upper_sprites_r),
.in_bitmap_display(in_bitmap_display),
.in_bitmap(in_bitmap_r),
.in_lower_sprites_display(in_lower_sprites_display),
.in_lower_sprites(in_lower_sprites_r),
.in_tilemap_display(in_tilemap_display),
.in_tilemap(in_tilemap_r),
.in_background(in_background_r),
.out_pix(_w_RED_pix),
.out_done(_w_RED_done),
.in_run(_RED_run),
.reset(reset),
.clock(clock)
);
M_expandcolour GREEN (
.in_terminal_display(in_terminal_display),
.in_terminal(in_terminal_g),
.in_character_map_display(in_character_map_display),
.in_character_map(in_character_map_g),
.in_upper_sprites_display(in_upper_sprites_display),
.in_upper_sprites(in_upper_sprites_g),
.in_bitmap_display(in_bitmap_display),
.in_bitmap(in_bitmap_g),
.in_lower_sprites_display(in_lower_sprites_display),
.in_lower_sprites(in_lower_sprites_g),
.in_tilemap_display(in_tilemap_display),
.in_tilemap(in_tilemap_g),
.in_background(in_background_g),
.out_pix(_w_GREEN_pix),
.out_done(_w_GREEN_done),
.in_run(_GREEN_run),
.reset(reset),
.clock(clock)
);
M_expandcolour BLUE (
.in_terminal_display(in_terminal_display),
.in_terminal(in_terminal_b),
.in_character_map_display(in_character_map_display),
.in_character_map(in_character_map_b),
.in_upper_sprites_display(in_upper_sprites_display),
.in_upper_sprites(in_upper_sprites_b),
.in_bitmap_display(in_bitmap_display),
.in_bitmap(in_bitmap_b),
.in_lower_sprites_display(in_lower_sprites_display),
.in_lower_sprites(in_lower_sprites_b),
.in_tilemap_display(in_tilemap_display),
.in_tilemap(in_tilemap_b),
.in_background(in_background_b),
.out_pix(_w_BLUE_pix),
.out_done(_w_BLUE_done),
.in_run(_BLUE_run),
.reset(reset),
.clock(clock)
);



always @* begin
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_index = _q_index;
_RED_run = 1;
_GREEN_run = 1;
_BLUE_run = 1;
// _always_pre
_d_pix_red = 0;
_d_pix_green = 0;
_d_pix_blue = 0;
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_pix_active) begin
// __block_5
// __block_7
_d_pix_red = _w_RED_pix;
_d_pix_green = _w_GREEN_pix;
_d_pix_blue = _w_BLUE_pix;
// __block_8
end else begin
// __block_6
end
// __block_9
// __block_10
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of multiplex_display
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_expandcolour (
in_terminal_display,
in_terminal,
in_character_map_display,
in_character_map,
in_upper_sprites_display,
in_upper_sprites,
in_bitmap_display,
in_bitmap,
in_lower_sprites_display,
in_lower_sprites,
in_tilemap_display,
in_tilemap,
in_background,
out_pix,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [0:0] in_terminal_display;
input  [1:0] in_terminal;
input  [0:0] in_character_map_display;
input  [1:0] in_character_map;
input  [0:0] in_upper_sprites_display;
input  [1:0] in_upper_sprites;
input  [0:0] in_bitmap_display;
input  [1:0] in_bitmap;
input  [0:0] in_lower_sprites_display;
input  [1:0] in_lower_sprites;
input  [0:0] in_tilemap_display;
input  [1:0] in_tilemap;
input  [1:0] in_background;
output  [7:0] out_pix;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [7:0] _d_pix,_q_pix;
reg  [1:0] _d_index,_q_index;
assign out_pix = _d_pix;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_pix <= _d_pix;
_q_index <= _d_index;
  end
end




always @* begin
_d_pix = _q_pix;
_d_index = _q_index;
// _always_pre
_d_pix = (in_terminal_display)?{{4{in_terminal}}}:(in_character_map_display)?{{4{in_character_map}}}:(in_upper_sprites_display)?{{4{in_upper_sprites}}}:(in_bitmap_display)?{{4{in_bitmap}}}:(in_lower_sprites_display)?{{4{in_lower_sprites}}}:(in_tilemap_display)?{{4{in_tilemap}}}:{{4{in_background}}};
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
// __block_5
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of expandcolour
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_pulse1hz (
in_resetCounter,
out_counter1hz,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [0:0] in_resetCounter;
output  [15:0] out_counter1hz;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [25:0] _d_counter50mhz;
reg  [25:0] _q_counter50mhz;
reg  [15:0] _d_counter1hz,_q_counter1hz;
reg  [1:0] _d_index,_q_index;
assign out_counter1hz = _q_counter1hz;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_counter50mhz <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_counter50mhz <= _d_counter50mhz;
_q_counter1hz <= _d_counter1hz;
_q_index <= _d_index;
  end
end




always @* begin
_d_counter50mhz = _q_counter50mhz;
_d_counter1hz = _q_counter1hz;
_d_index = _q_index;
// _always_pre
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_counter50mhz = 0;
// --
_d_counter1hz = 0;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_resetCounter==1) begin
// __block_5
// __block_7
_d_counter1hz = 0;
_d_counter50mhz = 0;
// __block_8
end else begin
// __block_6
// __block_9
_d_counter1hz = (_q_counter50mhz==50000000)?_q_counter1hz+1:_q_counter1hz;
_d_counter50mhz = (_q_counter50mhz==50000000)?0:_q_counter50mhz+1;
// __block_10
end
// __block_11
// __block_12
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of pulse1hz
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_pulse1khz (
in_resetCount,
in_resetCounter,
out_counter1khz,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_resetCount;
input  [0:0] in_resetCounter;
output  [15:0] out_counter1khz;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [15:0] _d_counter50mhz;
reg  [15:0] _q_counter50mhz;
reg  [15:0] _d_counter1khz,_q_counter1khz;
reg  [1:0] _d_index,_q_index;
assign out_counter1khz = _q_counter1khz;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_counter50mhz <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_counter50mhz <= _d_counter50mhz;
_q_counter1khz <= _d_counter1khz;
_q_index <= _d_index;
  end
end




always @* begin
_d_counter50mhz = _q_counter50mhz;
_d_counter1khz = _q_counter1khz;
_d_index = _q_index;
// _always_pre
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_counter50mhz = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_resetCounter==1) begin
// __block_5
// __block_7
_d_counter1khz = in_resetCount;
_d_counter50mhz = 0;
// __block_8
end else begin
// __block_6
// __block_9
_d_counter1khz = (_q_counter1khz==0)?0:(_q_counter50mhz==50000)?_q_counter1khz-1:_q_counter1khz;
_d_counter50mhz = (_q_counter50mhz==50000)?0:_q_counter50mhz+1;
// __block_10
end
// __block_11
// __block_12
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of pulse1khz
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_random (
in_resetRandom,
out_g_noise_out,
out_u_noise_out,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [0:0] in_resetRandom;
output  [15:0] out_g_noise_out;
output  [15:0] out_u_noise_out;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
reg  [15:0] _t_temp_u_noise3;
reg  [15:0] _t_temp_u_noise2;
reg  [15:0] _t_temp_u_noise1;
reg  [15:0] _t_temp_u_noise0;

reg  [15:0] _d_rand_out;
reg  [15:0] _q_rand_out;
reg  [15:0] _d_rand_ff;
reg  [15:0] _q_rand_ff;
reg  [17:0] _d_rand_en_ff;
reg  [17:0] _q_rand_en_ff;
reg  [15:0] _d_temp_g_noise_nxt;
reg  [15:0] _q_temp_g_noise_nxt;
reg  [15:0] _d_g_noise_out,_q_g_noise_out;
reg  [15:0] _d_u_noise_out,_q_u_noise_out;
reg  [1:0] _d_index,_q_index;
assign out_g_noise_out = _q_g_noise_out;
assign out_u_noise_out = _q_u_noise_out;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_rand_out <= 0;
_q_rand_ff <= 24'b011000110111011010011101;
_q_rand_en_ff <= 24'b001100010011011101100101;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_rand_out <= _d_rand_out;
_q_rand_ff <= _d_rand_ff;
_q_rand_en_ff <= _d_rand_en_ff;
_q_temp_g_noise_nxt <= _d_temp_g_noise_nxt;
_q_g_noise_out <= _d_g_noise_out;
_q_u_noise_out <= _d_u_noise_out;
_q_index <= _d_index;
  end
end




always @* begin
_d_rand_out = _q_rand_out;
_d_rand_ff = _q_rand_ff;
_d_rand_en_ff = _q_rand_en_ff;
_d_temp_g_noise_nxt = _q_temp_g_noise_nxt;
_d_g_noise_out = _q_g_noise_out;
_d_u_noise_out = _q_u_noise_out;
_d_index = _q_index;
_t_temp_u_noise3 = 0;
_t_temp_u_noise2 = 0;
_t_temp_u_noise1 = 0;
_t_temp_u_noise0 = 0;
// _always_pre
_d_g_noise_out = (_q_rand_en_ff[17+:1])?_q_temp_g_noise_nxt:(_q_rand_en_ff[10+:1])?_q_rand_out:_q_g_noise_out;
_d_u_noise_out = (_q_rand_en_ff[17+:1])?_q_rand_out:_q_u_noise_out;
_d_rand_en_ff = {(_q_rand_en_ff[7+:1]^_q_rand_en_ff[0+:1]),_q_rand_en_ff[1+:17]};
_d_rand_ff = {(_q_rand_ff[5+:1]^_q_rand_ff[3+:1]^_q_rand_ff[2+:1]^_q_rand_ff[0+:1]),_q_rand_ff[1+:15]};
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_rand_out = 0;
_d_rand_ff = 24'b011000110111011010011101;
_d_rand_en_ff = 24'b001100010011011101100101;
_t_temp_u_noise3 = 0;
_t_temp_u_noise2 = 0;
_t_temp_u_noise1 = 0;
_t_temp_u_noise0 = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_resetRandom) begin
// __block_5
// __block_7
_d_rand_en_ff = 24'b001100010011011101100101;
_d_rand_ff = 24'b011000110111011010011101;
_d_rand_out = 0;
_t_temp_u_noise3 = 0;
_t_temp_u_noise2 = 0;
_t_temp_u_noise1 = 0;
_t_temp_u_noise0 = 0;
_d_g_noise_out = 0;
_d_u_noise_out = 0;
// __block_8
end else begin
// __block_6
// __block_9
_d_rand_out = _d_rand_ff;
_t_temp_u_noise3 = {_d_rand_out[15+:1],_d_rand_out[15+:1],_d_rand_out[2+:13]};
_t_temp_u_noise2 = _t_temp_u_noise3;
_t_temp_u_noise1 = _t_temp_u_noise2;
_t_temp_u_noise0 = _t_temp_u_noise1;
_d_temp_g_noise_nxt = $signed(_t_temp_u_noise3)+$signed(_t_temp_u_noise2)+$signed(_t_temp_u_noise1)+$signed(_t_temp_u_noise0)+(_d_rand_en_ff[9+:1]?$signed(_d_g_noise_out):0);
// __block_10
end
// __block_11
// __block_12
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of random
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_terminal_mem_characterGenerator8x8(
input                  [10:0] in_characterGenerator8x8_addr,
output reg  [7:0] out_characterGenerator8x8_rdata,
input                                   clock
);
reg  [7:0] buffer[2047:0];
always @(posedge clock) begin
   out_characterGenerator8x8_rdata <= buffer[in_characterGenerator8x8_addr];
end
initial begin
 buffer[0] = 8'h00;
 buffer[1] = 8'h00;
 buffer[2] = 8'h00;
 buffer[3] = 8'h00;
 buffer[4] = 8'h00;
 buffer[5] = 8'h00;
 buffer[6] = 8'h00;
 buffer[7] = 8'h00;
 buffer[8] = 8'h7e;
 buffer[9] = 8'h81;
 buffer[10] = 8'ha5;
 buffer[11] = 8'h81;
 buffer[12] = 8'hbd;
 buffer[13] = 8'h99;
 buffer[14] = 8'h81;
 buffer[15] = 8'h7e;
 buffer[16] = 8'h7e;
 buffer[17] = 8'hff;
 buffer[18] = 8'hdb;
 buffer[19] = 8'hff;
 buffer[20] = 8'hc3;
 buffer[21] = 8'he7;
 buffer[22] = 8'hff;
 buffer[23] = 8'h7e;
 buffer[24] = 8'h6c;
 buffer[25] = 8'hfe;
 buffer[26] = 8'hfe;
 buffer[27] = 8'hfe;
 buffer[28] = 8'h7c;
 buffer[29] = 8'h38;
 buffer[30] = 8'h10;
 buffer[31] = 8'h00;
 buffer[32] = 8'h10;
 buffer[33] = 8'h38;
 buffer[34] = 8'h7c;
 buffer[35] = 8'hfe;
 buffer[36] = 8'h7c;
 buffer[37] = 8'h38;
 buffer[38] = 8'h10;
 buffer[39] = 8'h00;
 buffer[40] = 8'h38;
 buffer[41] = 8'h7c;
 buffer[42] = 8'h38;
 buffer[43] = 8'hfe;
 buffer[44] = 8'hfe;
 buffer[45] = 8'h7c;
 buffer[46] = 8'h38;
 buffer[47] = 8'h7c;
 buffer[48] = 8'h10;
 buffer[49] = 8'h10;
 buffer[50] = 8'h38;
 buffer[51] = 8'h7c;
 buffer[52] = 8'hfe;
 buffer[53] = 8'h7c;
 buffer[54] = 8'h38;
 buffer[55] = 8'h7c;
 buffer[56] = 8'h00;
 buffer[57] = 8'h00;
 buffer[58] = 8'h18;
 buffer[59] = 8'h3c;
 buffer[60] = 8'h3c;
 buffer[61] = 8'h18;
 buffer[62] = 8'h00;
 buffer[63] = 8'h00;
 buffer[64] = 8'hff;
 buffer[65] = 8'hff;
 buffer[66] = 8'he7;
 buffer[67] = 8'hc3;
 buffer[68] = 8'hc3;
 buffer[69] = 8'he7;
 buffer[70] = 8'hff;
 buffer[71] = 8'hff;
 buffer[72] = 8'h00;
 buffer[73] = 8'h3c;
 buffer[74] = 8'h66;
 buffer[75] = 8'h42;
 buffer[76] = 8'h42;
 buffer[77] = 8'h66;
 buffer[78] = 8'h3c;
 buffer[79] = 8'h00;
 buffer[80] = 8'hff;
 buffer[81] = 8'hc3;
 buffer[82] = 8'h99;
 buffer[83] = 8'hbd;
 buffer[84] = 8'hbd;
 buffer[85] = 8'h99;
 buffer[86] = 8'hc3;
 buffer[87] = 8'hff;
 buffer[88] = 8'h0f;
 buffer[89] = 8'h07;
 buffer[90] = 8'h0f;
 buffer[91] = 8'h7d;
 buffer[92] = 8'hcc;
 buffer[93] = 8'hcc;
 buffer[94] = 8'hcc;
 buffer[95] = 8'h78;
 buffer[96] = 8'h3c;
 buffer[97] = 8'h66;
 buffer[98] = 8'h66;
 buffer[99] = 8'h66;
 buffer[100] = 8'h3c;
 buffer[101] = 8'h18;
 buffer[102] = 8'h7e;
 buffer[103] = 8'h18;
 buffer[104] = 8'h3f;
 buffer[105] = 8'h33;
 buffer[106] = 8'h3f;
 buffer[107] = 8'h30;
 buffer[108] = 8'h30;
 buffer[109] = 8'h70;
 buffer[110] = 8'hf0;
 buffer[111] = 8'he0;
 buffer[112] = 8'h7f;
 buffer[113] = 8'h63;
 buffer[114] = 8'h7f;
 buffer[115] = 8'h63;
 buffer[116] = 8'h63;
 buffer[117] = 8'h67;
 buffer[118] = 8'he6;
 buffer[119] = 8'hc0;
 buffer[120] = 8'h99;
 buffer[121] = 8'h5a;
 buffer[122] = 8'h3c;
 buffer[123] = 8'he7;
 buffer[124] = 8'he7;
 buffer[125] = 8'h3c;
 buffer[126] = 8'h5a;
 buffer[127] = 8'h99;
 buffer[128] = 8'h80;
 buffer[129] = 8'he0;
 buffer[130] = 8'hf8;
 buffer[131] = 8'hfe;
 buffer[132] = 8'hf8;
 buffer[133] = 8'he0;
 buffer[134] = 8'h80;
 buffer[135] = 8'h00;
 buffer[136] = 8'h02;
 buffer[137] = 8'h0e;
 buffer[138] = 8'h3e;
 buffer[139] = 8'hfe;
 buffer[140] = 8'h3e;
 buffer[141] = 8'h0e;
 buffer[142] = 8'h02;
 buffer[143] = 8'h00;
 buffer[144] = 8'h18;
 buffer[145] = 8'h3c;
 buffer[146] = 8'h7e;
 buffer[147] = 8'h18;
 buffer[148] = 8'h18;
 buffer[149] = 8'h7e;
 buffer[150] = 8'h3c;
 buffer[151] = 8'h18;
 buffer[152] = 8'h66;
 buffer[153] = 8'h66;
 buffer[154] = 8'h66;
 buffer[155] = 8'h66;
 buffer[156] = 8'h66;
 buffer[157] = 8'h00;
 buffer[158] = 8'h66;
 buffer[159] = 8'h00;
 buffer[160] = 8'h7f;
 buffer[161] = 8'hdb;
 buffer[162] = 8'hdb;
 buffer[163] = 8'h7b;
 buffer[164] = 8'h1b;
 buffer[165] = 8'h1b;
 buffer[166] = 8'h1b;
 buffer[167] = 8'h00;
 buffer[168] = 8'h3e;
 buffer[169] = 8'h63;
 buffer[170] = 8'h38;
 buffer[171] = 8'h6c;
 buffer[172] = 8'h6c;
 buffer[173] = 8'h38;
 buffer[174] = 8'hcc;
 buffer[175] = 8'h78;
 buffer[176] = 8'h00;
 buffer[177] = 8'h00;
 buffer[178] = 8'h00;
 buffer[179] = 8'h00;
 buffer[180] = 8'h7e;
 buffer[181] = 8'h7e;
 buffer[182] = 8'h7e;
 buffer[183] = 8'h00;
 buffer[184] = 8'h18;
 buffer[185] = 8'h3c;
 buffer[186] = 8'h7e;
 buffer[187] = 8'h18;
 buffer[188] = 8'h7e;
 buffer[189] = 8'h3c;
 buffer[190] = 8'h18;
 buffer[191] = 8'hff;
 buffer[192] = 8'h18;
 buffer[193] = 8'h3c;
 buffer[194] = 8'h7e;
 buffer[195] = 8'h18;
 buffer[196] = 8'h18;
 buffer[197] = 8'h18;
 buffer[198] = 8'h18;
 buffer[199] = 8'h00;
 buffer[200] = 8'h18;
 buffer[201] = 8'h18;
 buffer[202] = 8'h18;
 buffer[203] = 8'h18;
 buffer[204] = 8'h7e;
 buffer[205] = 8'h3c;
 buffer[206] = 8'h18;
 buffer[207] = 8'h00;
 buffer[208] = 8'h00;
 buffer[209] = 8'h18;
 buffer[210] = 8'h0c;
 buffer[211] = 8'hfe;
 buffer[212] = 8'h0c;
 buffer[213] = 8'h18;
 buffer[214] = 8'h00;
 buffer[215] = 8'h00;
 buffer[216] = 8'h00;
 buffer[217] = 8'h30;
 buffer[218] = 8'h60;
 buffer[219] = 8'hfe;
 buffer[220] = 8'h60;
 buffer[221] = 8'h30;
 buffer[222] = 8'h00;
 buffer[223] = 8'h00;
 buffer[224] = 8'h00;
 buffer[225] = 8'h00;
 buffer[226] = 8'hc0;
 buffer[227] = 8'hc0;
 buffer[228] = 8'hc0;
 buffer[229] = 8'hfe;
 buffer[230] = 8'h00;
 buffer[231] = 8'h00;
 buffer[232] = 8'h00;
 buffer[233] = 8'h24;
 buffer[234] = 8'h66;
 buffer[235] = 8'hff;
 buffer[236] = 8'h66;
 buffer[237] = 8'h24;
 buffer[238] = 8'h00;
 buffer[239] = 8'h00;
 buffer[240] = 8'h00;
 buffer[241] = 8'h18;
 buffer[242] = 8'h3c;
 buffer[243] = 8'h7e;
 buffer[244] = 8'hff;
 buffer[245] = 8'hff;
 buffer[246] = 8'h00;
 buffer[247] = 8'h00;
 buffer[248] = 8'h00;
 buffer[249] = 8'hff;
 buffer[250] = 8'hff;
 buffer[251] = 8'h7e;
 buffer[252] = 8'h3c;
 buffer[253] = 8'h18;
 buffer[254] = 8'h00;
 buffer[255] = 8'h00;
 buffer[256] = 8'h00;
 buffer[257] = 8'h00;
 buffer[258] = 8'h00;
 buffer[259] = 8'h00;
 buffer[260] = 8'h00;
 buffer[261] = 8'h00;
 buffer[262] = 8'h00;
 buffer[263] = 8'h00;
 buffer[264] = 8'h30;
 buffer[265] = 8'h78;
 buffer[266] = 8'h78;
 buffer[267] = 8'h30;
 buffer[268] = 8'h30;
 buffer[269] = 8'h00;
 buffer[270] = 8'h30;
 buffer[271] = 8'h00;
 buffer[272] = 8'h6c;
 buffer[273] = 8'h6c;
 buffer[274] = 8'h6c;
 buffer[275] = 8'h00;
 buffer[276] = 8'h00;
 buffer[277] = 8'h00;
 buffer[278] = 8'h00;
 buffer[279] = 8'h00;
 buffer[280] = 8'h6c;
 buffer[281] = 8'h6c;
 buffer[282] = 8'hfe;
 buffer[283] = 8'h6c;
 buffer[284] = 8'hfe;
 buffer[285] = 8'h6c;
 buffer[286] = 8'h6c;
 buffer[287] = 8'h00;
 buffer[288] = 8'h30;
 buffer[289] = 8'h7c;
 buffer[290] = 8'hc0;
 buffer[291] = 8'h78;
 buffer[292] = 8'h0c;
 buffer[293] = 8'hf8;
 buffer[294] = 8'h30;
 buffer[295] = 8'h00;
 buffer[296] = 8'h00;
 buffer[297] = 8'hc6;
 buffer[298] = 8'hcc;
 buffer[299] = 8'h18;
 buffer[300] = 8'h30;
 buffer[301] = 8'h66;
 buffer[302] = 8'hc6;
 buffer[303] = 8'h00;
 buffer[304] = 8'h38;
 buffer[305] = 8'h6c;
 buffer[306] = 8'h38;
 buffer[307] = 8'h76;
 buffer[308] = 8'hdc;
 buffer[309] = 8'hcc;
 buffer[310] = 8'h76;
 buffer[311] = 8'h00;
 buffer[312] = 8'h60;
 buffer[313] = 8'h60;
 buffer[314] = 8'hc0;
 buffer[315] = 8'h00;
 buffer[316] = 8'h00;
 buffer[317] = 8'h00;
 buffer[318] = 8'h00;
 buffer[319] = 8'h00;
 buffer[320] = 8'h18;
 buffer[321] = 8'h30;
 buffer[322] = 8'h60;
 buffer[323] = 8'h60;
 buffer[324] = 8'h60;
 buffer[325] = 8'h30;
 buffer[326] = 8'h18;
 buffer[327] = 8'h00;
 buffer[328] = 8'h60;
 buffer[329] = 8'h30;
 buffer[330] = 8'h18;
 buffer[331] = 8'h18;
 buffer[332] = 8'h18;
 buffer[333] = 8'h30;
 buffer[334] = 8'h60;
 buffer[335] = 8'h00;
 buffer[336] = 8'h00;
 buffer[337] = 8'h66;
 buffer[338] = 8'h3c;
 buffer[339] = 8'hff;
 buffer[340] = 8'h3c;
 buffer[341] = 8'h66;
 buffer[342] = 8'h00;
 buffer[343] = 8'h00;
 buffer[344] = 8'h00;
 buffer[345] = 8'h30;
 buffer[346] = 8'h30;
 buffer[347] = 8'hfc;
 buffer[348] = 8'h30;
 buffer[349] = 8'h30;
 buffer[350] = 8'h00;
 buffer[351] = 8'h00;
 buffer[352] = 8'h00;
 buffer[353] = 8'h00;
 buffer[354] = 8'h00;
 buffer[355] = 8'h00;
 buffer[356] = 8'h00;
 buffer[357] = 8'h30;
 buffer[358] = 8'h30;
 buffer[359] = 8'h60;
 buffer[360] = 8'h00;
 buffer[361] = 8'h00;
 buffer[362] = 8'h00;
 buffer[363] = 8'hfc;
 buffer[364] = 8'h00;
 buffer[365] = 8'h00;
 buffer[366] = 8'h00;
 buffer[367] = 8'h00;
 buffer[368] = 8'h00;
 buffer[369] = 8'h00;
 buffer[370] = 8'h00;
 buffer[371] = 8'h00;
 buffer[372] = 8'h00;
 buffer[373] = 8'h30;
 buffer[374] = 8'h30;
 buffer[375] = 8'h00;
 buffer[376] = 8'h06;
 buffer[377] = 8'h0c;
 buffer[378] = 8'h18;
 buffer[379] = 8'h30;
 buffer[380] = 8'h60;
 buffer[381] = 8'hc0;
 buffer[382] = 8'h80;
 buffer[383] = 8'h00;
 buffer[384] = 8'h7c;
 buffer[385] = 8'hc6;
 buffer[386] = 8'hce;
 buffer[387] = 8'hde;
 buffer[388] = 8'hf6;
 buffer[389] = 8'he6;
 buffer[390] = 8'h7c;
 buffer[391] = 8'h00;
 buffer[392] = 8'h30;
 buffer[393] = 8'h70;
 buffer[394] = 8'h30;
 buffer[395] = 8'h30;
 buffer[396] = 8'h30;
 buffer[397] = 8'h30;
 buffer[398] = 8'hfc;
 buffer[399] = 8'h00;
 buffer[400] = 8'h78;
 buffer[401] = 8'hcc;
 buffer[402] = 8'h0c;
 buffer[403] = 8'h38;
 buffer[404] = 8'h60;
 buffer[405] = 8'hcc;
 buffer[406] = 8'hfc;
 buffer[407] = 8'h00;
 buffer[408] = 8'h78;
 buffer[409] = 8'hcc;
 buffer[410] = 8'h0c;
 buffer[411] = 8'h38;
 buffer[412] = 8'h0c;
 buffer[413] = 8'hcc;
 buffer[414] = 8'h78;
 buffer[415] = 8'h00;
 buffer[416] = 8'h1c;
 buffer[417] = 8'h3c;
 buffer[418] = 8'h6c;
 buffer[419] = 8'hcc;
 buffer[420] = 8'hfe;
 buffer[421] = 8'h0c;
 buffer[422] = 8'h1e;
 buffer[423] = 8'h00;
 buffer[424] = 8'hfc;
 buffer[425] = 8'hc0;
 buffer[426] = 8'hf8;
 buffer[427] = 8'h0c;
 buffer[428] = 8'h0c;
 buffer[429] = 8'hcc;
 buffer[430] = 8'h78;
 buffer[431] = 8'h00;
 buffer[432] = 8'h38;
 buffer[433] = 8'h60;
 buffer[434] = 8'hc0;
 buffer[435] = 8'hf8;
 buffer[436] = 8'hcc;
 buffer[437] = 8'hcc;
 buffer[438] = 8'h78;
 buffer[439] = 8'h00;
 buffer[440] = 8'hfc;
 buffer[441] = 8'hcc;
 buffer[442] = 8'h0c;
 buffer[443] = 8'h18;
 buffer[444] = 8'h30;
 buffer[445] = 8'h30;
 buffer[446] = 8'h30;
 buffer[447] = 8'h00;
 buffer[448] = 8'h78;
 buffer[449] = 8'hcc;
 buffer[450] = 8'hcc;
 buffer[451] = 8'h78;
 buffer[452] = 8'hcc;
 buffer[453] = 8'hcc;
 buffer[454] = 8'h78;
 buffer[455] = 8'h00;
 buffer[456] = 8'h78;
 buffer[457] = 8'hcc;
 buffer[458] = 8'hcc;
 buffer[459] = 8'h7c;
 buffer[460] = 8'h0c;
 buffer[461] = 8'h18;
 buffer[462] = 8'h70;
 buffer[463] = 8'h00;
 buffer[464] = 8'h00;
 buffer[465] = 8'h30;
 buffer[466] = 8'h30;
 buffer[467] = 8'h00;
 buffer[468] = 8'h00;
 buffer[469] = 8'h30;
 buffer[470] = 8'h30;
 buffer[471] = 8'h00;
 buffer[472] = 8'h00;
 buffer[473] = 8'h30;
 buffer[474] = 8'h30;
 buffer[475] = 8'h00;
 buffer[476] = 8'h00;
 buffer[477] = 8'h30;
 buffer[478] = 8'h30;
 buffer[479] = 8'h60;
 buffer[480] = 8'h18;
 buffer[481] = 8'h30;
 buffer[482] = 8'h60;
 buffer[483] = 8'hc0;
 buffer[484] = 8'h60;
 buffer[485] = 8'h30;
 buffer[486] = 8'h18;
 buffer[487] = 8'h00;
 buffer[488] = 8'h00;
 buffer[489] = 8'h00;
 buffer[490] = 8'hfc;
 buffer[491] = 8'h00;
 buffer[492] = 8'h00;
 buffer[493] = 8'hfc;
 buffer[494] = 8'h00;
 buffer[495] = 8'h00;
 buffer[496] = 8'h60;
 buffer[497] = 8'h30;
 buffer[498] = 8'h18;
 buffer[499] = 8'h0c;
 buffer[500] = 8'h18;
 buffer[501] = 8'h30;
 buffer[502] = 8'h60;
 buffer[503] = 8'h00;
 buffer[504] = 8'h78;
 buffer[505] = 8'hcc;
 buffer[506] = 8'h0c;
 buffer[507] = 8'h18;
 buffer[508] = 8'h30;
 buffer[509] = 8'h00;
 buffer[510] = 8'h30;
 buffer[511] = 8'h00;
 buffer[512] = 8'h7c;
 buffer[513] = 8'hc6;
 buffer[514] = 8'hde;
 buffer[515] = 8'hde;
 buffer[516] = 8'hde;
 buffer[517] = 8'hc0;
 buffer[518] = 8'h78;
 buffer[519] = 8'h00;
 buffer[520] = 8'h30;
 buffer[521] = 8'h78;
 buffer[522] = 8'hcc;
 buffer[523] = 8'hcc;
 buffer[524] = 8'hfc;
 buffer[525] = 8'hcc;
 buffer[526] = 8'hcc;
 buffer[527] = 8'h00;
 buffer[528] = 8'hfc;
 buffer[529] = 8'h66;
 buffer[530] = 8'h66;
 buffer[531] = 8'h7c;
 buffer[532] = 8'h66;
 buffer[533] = 8'h66;
 buffer[534] = 8'hfc;
 buffer[535] = 8'h00;
 buffer[536] = 8'h3c;
 buffer[537] = 8'h66;
 buffer[538] = 8'hc0;
 buffer[539] = 8'hc0;
 buffer[540] = 8'hc0;
 buffer[541] = 8'h66;
 buffer[542] = 8'h3c;
 buffer[543] = 8'h00;
 buffer[544] = 8'hf8;
 buffer[545] = 8'h6c;
 buffer[546] = 8'h66;
 buffer[547] = 8'h66;
 buffer[548] = 8'h66;
 buffer[549] = 8'h6c;
 buffer[550] = 8'hf8;
 buffer[551] = 8'h00;
 buffer[552] = 8'hfe;
 buffer[553] = 8'h62;
 buffer[554] = 8'h68;
 buffer[555] = 8'h78;
 buffer[556] = 8'h68;
 buffer[557] = 8'h62;
 buffer[558] = 8'hfe;
 buffer[559] = 8'h00;
 buffer[560] = 8'hfe;
 buffer[561] = 8'h62;
 buffer[562] = 8'h68;
 buffer[563] = 8'h78;
 buffer[564] = 8'h68;
 buffer[565] = 8'h60;
 buffer[566] = 8'hf0;
 buffer[567] = 8'h00;
 buffer[568] = 8'h3c;
 buffer[569] = 8'h66;
 buffer[570] = 8'hc0;
 buffer[571] = 8'hc0;
 buffer[572] = 8'hce;
 buffer[573] = 8'h66;
 buffer[574] = 8'h3e;
 buffer[575] = 8'h00;
 buffer[576] = 8'hcc;
 buffer[577] = 8'hcc;
 buffer[578] = 8'hcc;
 buffer[579] = 8'hfc;
 buffer[580] = 8'hcc;
 buffer[581] = 8'hcc;
 buffer[582] = 8'hcc;
 buffer[583] = 8'h00;
 buffer[584] = 8'h78;
 buffer[585] = 8'h30;
 buffer[586] = 8'h30;
 buffer[587] = 8'h30;
 buffer[588] = 8'h30;
 buffer[589] = 8'h30;
 buffer[590] = 8'h78;
 buffer[591] = 8'h00;
 buffer[592] = 8'h1e;
 buffer[593] = 8'h0c;
 buffer[594] = 8'h0c;
 buffer[595] = 8'h0c;
 buffer[596] = 8'hcc;
 buffer[597] = 8'hcc;
 buffer[598] = 8'h78;
 buffer[599] = 8'h00;
 buffer[600] = 8'he6;
 buffer[601] = 8'h66;
 buffer[602] = 8'h6c;
 buffer[603] = 8'h78;
 buffer[604] = 8'h6c;
 buffer[605] = 8'h66;
 buffer[606] = 8'he6;
 buffer[607] = 8'h00;
 buffer[608] = 8'hf0;
 buffer[609] = 8'h60;
 buffer[610] = 8'h60;
 buffer[611] = 8'h60;
 buffer[612] = 8'h62;
 buffer[613] = 8'h66;
 buffer[614] = 8'hfe;
 buffer[615] = 8'h00;
 buffer[616] = 8'hc6;
 buffer[617] = 8'hee;
 buffer[618] = 8'hfe;
 buffer[619] = 8'hfe;
 buffer[620] = 8'hd6;
 buffer[621] = 8'hc6;
 buffer[622] = 8'hc6;
 buffer[623] = 8'h00;
 buffer[624] = 8'hc6;
 buffer[625] = 8'he6;
 buffer[626] = 8'hf6;
 buffer[627] = 8'hde;
 buffer[628] = 8'hce;
 buffer[629] = 8'hc6;
 buffer[630] = 8'hc6;
 buffer[631] = 8'h00;
 buffer[632] = 8'h38;
 buffer[633] = 8'h6c;
 buffer[634] = 8'hc6;
 buffer[635] = 8'hc6;
 buffer[636] = 8'hc6;
 buffer[637] = 8'h6c;
 buffer[638] = 8'h38;
 buffer[639] = 8'h00;
 buffer[640] = 8'hfc;
 buffer[641] = 8'h66;
 buffer[642] = 8'h66;
 buffer[643] = 8'h7c;
 buffer[644] = 8'h60;
 buffer[645] = 8'h60;
 buffer[646] = 8'hf0;
 buffer[647] = 8'h00;
 buffer[648] = 8'h78;
 buffer[649] = 8'hcc;
 buffer[650] = 8'hcc;
 buffer[651] = 8'hcc;
 buffer[652] = 8'hdc;
 buffer[653] = 8'h78;
 buffer[654] = 8'h1c;
 buffer[655] = 8'h00;
 buffer[656] = 8'hfc;
 buffer[657] = 8'h66;
 buffer[658] = 8'h66;
 buffer[659] = 8'h7c;
 buffer[660] = 8'h6c;
 buffer[661] = 8'h66;
 buffer[662] = 8'he6;
 buffer[663] = 8'h00;
 buffer[664] = 8'h78;
 buffer[665] = 8'hcc;
 buffer[666] = 8'he0;
 buffer[667] = 8'h70;
 buffer[668] = 8'h1c;
 buffer[669] = 8'hcc;
 buffer[670] = 8'h78;
 buffer[671] = 8'h00;
 buffer[672] = 8'hfc;
 buffer[673] = 8'hb4;
 buffer[674] = 8'h30;
 buffer[675] = 8'h30;
 buffer[676] = 8'h30;
 buffer[677] = 8'h30;
 buffer[678] = 8'h78;
 buffer[679] = 8'h00;
 buffer[680] = 8'hcc;
 buffer[681] = 8'hcc;
 buffer[682] = 8'hcc;
 buffer[683] = 8'hcc;
 buffer[684] = 8'hcc;
 buffer[685] = 8'hcc;
 buffer[686] = 8'hfc;
 buffer[687] = 8'h00;
 buffer[688] = 8'hcc;
 buffer[689] = 8'hcc;
 buffer[690] = 8'hcc;
 buffer[691] = 8'hcc;
 buffer[692] = 8'hcc;
 buffer[693] = 8'h78;
 buffer[694] = 8'h30;
 buffer[695] = 8'h00;
 buffer[696] = 8'hc6;
 buffer[697] = 8'hc6;
 buffer[698] = 8'hc6;
 buffer[699] = 8'hd6;
 buffer[700] = 8'hfe;
 buffer[701] = 8'hee;
 buffer[702] = 8'hc6;
 buffer[703] = 8'h00;
 buffer[704] = 8'hc6;
 buffer[705] = 8'hc6;
 buffer[706] = 8'h6c;
 buffer[707] = 8'h38;
 buffer[708] = 8'h38;
 buffer[709] = 8'h6c;
 buffer[710] = 8'hc6;
 buffer[711] = 8'h00;
 buffer[712] = 8'hcc;
 buffer[713] = 8'hcc;
 buffer[714] = 8'hcc;
 buffer[715] = 8'h78;
 buffer[716] = 8'h30;
 buffer[717] = 8'h30;
 buffer[718] = 8'h78;
 buffer[719] = 8'h00;
 buffer[720] = 8'hfe;
 buffer[721] = 8'hc6;
 buffer[722] = 8'h8c;
 buffer[723] = 8'h18;
 buffer[724] = 8'h32;
 buffer[725] = 8'h66;
 buffer[726] = 8'hfe;
 buffer[727] = 8'h00;
 buffer[728] = 8'h78;
 buffer[729] = 8'h60;
 buffer[730] = 8'h60;
 buffer[731] = 8'h60;
 buffer[732] = 8'h60;
 buffer[733] = 8'h60;
 buffer[734] = 8'h78;
 buffer[735] = 8'h00;
 buffer[736] = 8'hc0;
 buffer[737] = 8'h60;
 buffer[738] = 8'h30;
 buffer[739] = 8'h18;
 buffer[740] = 8'h0c;
 buffer[741] = 8'h06;
 buffer[742] = 8'h02;
 buffer[743] = 8'h00;
 buffer[744] = 8'h78;
 buffer[745] = 8'h18;
 buffer[746] = 8'h18;
 buffer[747] = 8'h18;
 buffer[748] = 8'h18;
 buffer[749] = 8'h18;
 buffer[750] = 8'h78;
 buffer[751] = 8'h00;
 buffer[752] = 8'h10;
 buffer[753] = 8'h38;
 buffer[754] = 8'h6c;
 buffer[755] = 8'hc6;
 buffer[756] = 8'h00;
 buffer[757] = 8'h00;
 buffer[758] = 8'h00;
 buffer[759] = 8'h00;
 buffer[760] = 8'h00;
 buffer[761] = 8'h00;
 buffer[762] = 8'h00;
 buffer[763] = 8'h00;
 buffer[764] = 8'h00;
 buffer[765] = 8'h00;
 buffer[766] = 8'h00;
 buffer[767] = 8'hff;
 buffer[768] = 8'h30;
 buffer[769] = 8'h30;
 buffer[770] = 8'h18;
 buffer[771] = 8'h00;
 buffer[772] = 8'h00;
 buffer[773] = 8'h00;
 buffer[774] = 8'h00;
 buffer[775] = 8'h00;
 buffer[776] = 8'h00;
 buffer[777] = 8'h00;
 buffer[778] = 8'h78;
 buffer[779] = 8'h0c;
 buffer[780] = 8'h7c;
 buffer[781] = 8'hcc;
 buffer[782] = 8'h76;
 buffer[783] = 8'h00;
 buffer[784] = 8'he0;
 buffer[785] = 8'h60;
 buffer[786] = 8'h60;
 buffer[787] = 8'h7c;
 buffer[788] = 8'h66;
 buffer[789] = 8'h66;
 buffer[790] = 8'hdc;
 buffer[791] = 8'h00;
 buffer[792] = 8'h00;
 buffer[793] = 8'h00;
 buffer[794] = 8'h78;
 buffer[795] = 8'hcc;
 buffer[796] = 8'hc0;
 buffer[797] = 8'hcc;
 buffer[798] = 8'h78;
 buffer[799] = 8'h00;
 buffer[800] = 8'h1c;
 buffer[801] = 8'h0c;
 buffer[802] = 8'h0c;
 buffer[803] = 8'h7c;
 buffer[804] = 8'hcc;
 buffer[805] = 8'hcc;
 buffer[806] = 8'h76;
 buffer[807] = 8'h00;
 buffer[808] = 8'h00;
 buffer[809] = 8'h00;
 buffer[810] = 8'h78;
 buffer[811] = 8'hcc;
 buffer[812] = 8'hfc;
 buffer[813] = 8'hc0;
 buffer[814] = 8'h78;
 buffer[815] = 8'h00;
 buffer[816] = 8'h38;
 buffer[817] = 8'h6c;
 buffer[818] = 8'h60;
 buffer[819] = 8'hf0;
 buffer[820] = 8'h60;
 buffer[821] = 8'h60;
 buffer[822] = 8'hf0;
 buffer[823] = 8'h00;
 buffer[824] = 8'h00;
 buffer[825] = 8'h00;
 buffer[826] = 8'h76;
 buffer[827] = 8'hcc;
 buffer[828] = 8'hcc;
 buffer[829] = 8'h7c;
 buffer[830] = 8'h0c;
 buffer[831] = 8'hf8;
 buffer[832] = 8'he0;
 buffer[833] = 8'h60;
 buffer[834] = 8'h6c;
 buffer[835] = 8'h76;
 buffer[836] = 8'h66;
 buffer[837] = 8'h66;
 buffer[838] = 8'he6;
 buffer[839] = 8'h00;
 buffer[840] = 8'h30;
 buffer[841] = 8'h00;
 buffer[842] = 8'h70;
 buffer[843] = 8'h30;
 buffer[844] = 8'h30;
 buffer[845] = 8'h30;
 buffer[846] = 8'h78;
 buffer[847] = 8'h00;
 buffer[848] = 8'h0c;
 buffer[849] = 8'h00;
 buffer[850] = 8'h0c;
 buffer[851] = 8'h0c;
 buffer[852] = 8'h0c;
 buffer[853] = 8'hcc;
 buffer[854] = 8'hcc;
 buffer[855] = 8'h78;
 buffer[856] = 8'he0;
 buffer[857] = 8'h60;
 buffer[858] = 8'h66;
 buffer[859] = 8'h6c;
 buffer[860] = 8'h78;
 buffer[861] = 8'h6c;
 buffer[862] = 8'he6;
 buffer[863] = 8'h00;
 buffer[864] = 8'h70;
 buffer[865] = 8'h30;
 buffer[866] = 8'h30;
 buffer[867] = 8'h30;
 buffer[868] = 8'h30;
 buffer[869] = 8'h30;
 buffer[870] = 8'h78;
 buffer[871] = 8'h00;
 buffer[872] = 8'h00;
 buffer[873] = 8'h00;
 buffer[874] = 8'hcc;
 buffer[875] = 8'hfe;
 buffer[876] = 8'hfe;
 buffer[877] = 8'hd6;
 buffer[878] = 8'hc6;
 buffer[879] = 8'h00;
 buffer[880] = 8'h00;
 buffer[881] = 8'h00;
 buffer[882] = 8'hf8;
 buffer[883] = 8'hcc;
 buffer[884] = 8'hcc;
 buffer[885] = 8'hcc;
 buffer[886] = 8'hcc;
 buffer[887] = 8'h00;
 buffer[888] = 8'h00;
 buffer[889] = 8'h00;
 buffer[890] = 8'h78;
 buffer[891] = 8'hcc;
 buffer[892] = 8'hcc;
 buffer[893] = 8'hcc;
 buffer[894] = 8'h78;
 buffer[895] = 8'h00;
 buffer[896] = 8'h00;
 buffer[897] = 8'h00;
 buffer[898] = 8'hdc;
 buffer[899] = 8'h66;
 buffer[900] = 8'h66;
 buffer[901] = 8'h7c;
 buffer[902] = 8'h60;
 buffer[903] = 8'hf0;
 buffer[904] = 8'h00;
 buffer[905] = 8'h00;
 buffer[906] = 8'h76;
 buffer[907] = 8'hcc;
 buffer[908] = 8'hcc;
 buffer[909] = 8'h7c;
 buffer[910] = 8'h0c;
 buffer[911] = 8'h1e;
 buffer[912] = 8'h00;
 buffer[913] = 8'h00;
 buffer[914] = 8'hdc;
 buffer[915] = 8'h76;
 buffer[916] = 8'h66;
 buffer[917] = 8'h60;
 buffer[918] = 8'hf0;
 buffer[919] = 8'h00;
 buffer[920] = 8'h00;
 buffer[921] = 8'h00;
 buffer[922] = 8'h7c;
 buffer[923] = 8'hc0;
 buffer[924] = 8'h78;
 buffer[925] = 8'h0c;
 buffer[926] = 8'hf8;
 buffer[927] = 8'h00;
 buffer[928] = 8'h10;
 buffer[929] = 8'h30;
 buffer[930] = 8'h7c;
 buffer[931] = 8'h30;
 buffer[932] = 8'h30;
 buffer[933] = 8'h34;
 buffer[934] = 8'h18;
 buffer[935] = 8'h00;
 buffer[936] = 8'h00;
 buffer[937] = 8'h00;
 buffer[938] = 8'hcc;
 buffer[939] = 8'hcc;
 buffer[940] = 8'hcc;
 buffer[941] = 8'hcc;
 buffer[942] = 8'h76;
 buffer[943] = 8'h00;
 buffer[944] = 8'h00;
 buffer[945] = 8'h00;
 buffer[946] = 8'hcc;
 buffer[947] = 8'hcc;
 buffer[948] = 8'hcc;
 buffer[949] = 8'h78;
 buffer[950] = 8'h30;
 buffer[951] = 8'h00;
 buffer[952] = 8'h00;
 buffer[953] = 8'h00;
 buffer[954] = 8'hc6;
 buffer[955] = 8'hd6;
 buffer[956] = 8'hfe;
 buffer[957] = 8'hfe;
 buffer[958] = 8'h6c;
 buffer[959] = 8'h00;
 buffer[960] = 8'h00;
 buffer[961] = 8'h00;
 buffer[962] = 8'hc6;
 buffer[963] = 8'h6c;
 buffer[964] = 8'h38;
 buffer[965] = 8'h6c;
 buffer[966] = 8'hc6;
 buffer[967] = 8'h00;
 buffer[968] = 8'h00;
 buffer[969] = 8'h00;
 buffer[970] = 8'hcc;
 buffer[971] = 8'hcc;
 buffer[972] = 8'hcc;
 buffer[973] = 8'h7c;
 buffer[974] = 8'h0c;
 buffer[975] = 8'hf8;
 buffer[976] = 8'h00;
 buffer[977] = 8'h00;
 buffer[978] = 8'hfc;
 buffer[979] = 8'h98;
 buffer[980] = 8'h30;
 buffer[981] = 8'h64;
 buffer[982] = 8'hfc;
 buffer[983] = 8'h00;
 buffer[984] = 8'h1c;
 buffer[985] = 8'h30;
 buffer[986] = 8'h30;
 buffer[987] = 8'he0;
 buffer[988] = 8'h30;
 buffer[989] = 8'h30;
 buffer[990] = 8'h1c;
 buffer[991] = 8'h00;
 buffer[992] = 8'h18;
 buffer[993] = 8'h18;
 buffer[994] = 8'h18;
 buffer[995] = 8'h00;
 buffer[996] = 8'h18;
 buffer[997] = 8'h18;
 buffer[998] = 8'h18;
 buffer[999] = 8'h00;
 buffer[1000] = 8'he0;
 buffer[1001] = 8'h30;
 buffer[1002] = 8'h30;
 buffer[1003] = 8'h1c;
 buffer[1004] = 8'h30;
 buffer[1005] = 8'h30;
 buffer[1006] = 8'he0;
 buffer[1007] = 8'h00;
 buffer[1008] = 8'h76;
 buffer[1009] = 8'hdc;
 buffer[1010] = 8'h00;
 buffer[1011] = 8'h00;
 buffer[1012] = 8'h00;
 buffer[1013] = 8'h00;
 buffer[1014] = 8'h00;
 buffer[1015] = 8'h00;
 buffer[1016] = 8'h00;
 buffer[1017] = 8'h10;
 buffer[1018] = 8'h38;
 buffer[1019] = 8'h6c;
 buffer[1020] = 8'hc6;
 buffer[1021] = 8'hc6;
 buffer[1022] = 8'hfe;
 buffer[1023] = 8'h00;
 buffer[1024] = 8'h78;
 buffer[1025] = 8'hcc;
 buffer[1026] = 8'hc0;
 buffer[1027] = 8'hcc;
 buffer[1028] = 8'h78;
 buffer[1029] = 8'h18;
 buffer[1030] = 8'h0c;
 buffer[1031] = 8'h78;
 buffer[1032] = 8'h00;
 buffer[1033] = 8'hcc;
 buffer[1034] = 8'h00;
 buffer[1035] = 8'hcc;
 buffer[1036] = 8'hcc;
 buffer[1037] = 8'hcc;
 buffer[1038] = 8'h7e;
 buffer[1039] = 8'h00;
 buffer[1040] = 8'h1c;
 buffer[1041] = 8'h00;
 buffer[1042] = 8'h78;
 buffer[1043] = 8'hcc;
 buffer[1044] = 8'hfc;
 buffer[1045] = 8'hc0;
 buffer[1046] = 8'h78;
 buffer[1047] = 8'h00;
 buffer[1048] = 8'h7e;
 buffer[1049] = 8'hc3;
 buffer[1050] = 8'h3c;
 buffer[1051] = 8'h06;
 buffer[1052] = 8'h3e;
 buffer[1053] = 8'h66;
 buffer[1054] = 8'h3f;
 buffer[1055] = 8'h00;
 buffer[1056] = 8'hcc;
 buffer[1057] = 8'h00;
 buffer[1058] = 8'h78;
 buffer[1059] = 8'h0c;
 buffer[1060] = 8'h7c;
 buffer[1061] = 8'hcc;
 buffer[1062] = 8'h7e;
 buffer[1063] = 8'h00;
 buffer[1064] = 8'he0;
 buffer[1065] = 8'h00;
 buffer[1066] = 8'h78;
 buffer[1067] = 8'h0c;
 buffer[1068] = 8'h7c;
 buffer[1069] = 8'hcc;
 buffer[1070] = 8'h7e;
 buffer[1071] = 8'h00;
 buffer[1072] = 8'h30;
 buffer[1073] = 8'h30;
 buffer[1074] = 8'h78;
 buffer[1075] = 8'h0c;
 buffer[1076] = 8'h7c;
 buffer[1077] = 8'hcc;
 buffer[1078] = 8'h7e;
 buffer[1079] = 8'h00;
 buffer[1080] = 8'h00;
 buffer[1081] = 8'h00;
 buffer[1082] = 8'h78;
 buffer[1083] = 8'hc0;
 buffer[1084] = 8'hc0;
 buffer[1085] = 8'h78;
 buffer[1086] = 8'h0c;
 buffer[1087] = 8'h38;
 buffer[1088] = 8'h7e;
 buffer[1089] = 8'hc3;
 buffer[1090] = 8'h3c;
 buffer[1091] = 8'h66;
 buffer[1092] = 8'h7e;
 buffer[1093] = 8'h60;
 buffer[1094] = 8'h3c;
 buffer[1095] = 8'h00;
 buffer[1096] = 8'hcc;
 buffer[1097] = 8'h00;
 buffer[1098] = 8'h78;
 buffer[1099] = 8'hcc;
 buffer[1100] = 8'hfc;
 buffer[1101] = 8'hc0;
 buffer[1102] = 8'h78;
 buffer[1103] = 8'h00;
 buffer[1104] = 8'he0;
 buffer[1105] = 8'h00;
 buffer[1106] = 8'h78;
 buffer[1107] = 8'hcc;
 buffer[1108] = 8'hfc;
 buffer[1109] = 8'hc0;
 buffer[1110] = 8'h78;
 buffer[1111] = 8'h00;
 buffer[1112] = 8'hcc;
 buffer[1113] = 8'h00;
 buffer[1114] = 8'h70;
 buffer[1115] = 8'h30;
 buffer[1116] = 8'h30;
 buffer[1117] = 8'h30;
 buffer[1118] = 8'h78;
 buffer[1119] = 8'h00;
 buffer[1120] = 8'h7c;
 buffer[1121] = 8'hc6;
 buffer[1122] = 8'h38;
 buffer[1123] = 8'h18;
 buffer[1124] = 8'h18;
 buffer[1125] = 8'h18;
 buffer[1126] = 8'h3c;
 buffer[1127] = 8'h00;
 buffer[1128] = 8'he0;
 buffer[1129] = 8'h00;
 buffer[1130] = 8'h70;
 buffer[1131] = 8'h30;
 buffer[1132] = 8'h30;
 buffer[1133] = 8'h30;
 buffer[1134] = 8'h78;
 buffer[1135] = 8'h00;
 buffer[1136] = 8'hc6;
 buffer[1137] = 8'h38;
 buffer[1138] = 8'h6c;
 buffer[1139] = 8'hc6;
 buffer[1140] = 8'hfe;
 buffer[1141] = 8'hc6;
 buffer[1142] = 8'hc6;
 buffer[1143] = 8'h00;
 buffer[1144] = 8'h30;
 buffer[1145] = 8'h30;
 buffer[1146] = 8'h00;
 buffer[1147] = 8'h78;
 buffer[1148] = 8'hcc;
 buffer[1149] = 8'hfc;
 buffer[1150] = 8'hcc;
 buffer[1151] = 8'h00;
 buffer[1152] = 8'h1c;
 buffer[1153] = 8'h00;
 buffer[1154] = 8'hfc;
 buffer[1155] = 8'h60;
 buffer[1156] = 8'h78;
 buffer[1157] = 8'h60;
 buffer[1158] = 8'hfc;
 buffer[1159] = 8'h00;
 buffer[1160] = 8'h00;
 buffer[1161] = 8'h00;
 buffer[1162] = 8'h7f;
 buffer[1163] = 8'h0c;
 buffer[1164] = 8'h7f;
 buffer[1165] = 8'hcc;
 buffer[1166] = 8'h7f;
 buffer[1167] = 8'h00;
 buffer[1168] = 8'h3e;
 buffer[1169] = 8'h6c;
 buffer[1170] = 8'hcc;
 buffer[1171] = 8'hfe;
 buffer[1172] = 8'hcc;
 buffer[1173] = 8'hcc;
 buffer[1174] = 8'hce;
 buffer[1175] = 8'h00;
 buffer[1176] = 8'h78;
 buffer[1177] = 8'hcc;
 buffer[1178] = 8'h00;
 buffer[1179] = 8'h78;
 buffer[1180] = 8'hcc;
 buffer[1181] = 8'hcc;
 buffer[1182] = 8'h78;
 buffer[1183] = 8'h00;
 buffer[1184] = 8'h00;
 buffer[1185] = 8'hcc;
 buffer[1186] = 8'h00;
 buffer[1187] = 8'h78;
 buffer[1188] = 8'hcc;
 buffer[1189] = 8'hcc;
 buffer[1190] = 8'h78;
 buffer[1191] = 8'h00;
 buffer[1192] = 8'h00;
 buffer[1193] = 8'he0;
 buffer[1194] = 8'h00;
 buffer[1195] = 8'h78;
 buffer[1196] = 8'hcc;
 buffer[1197] = 8'hcc;
 buffer[1198] = 8'h78;
 buffer[1199] = 8'h00;
 buffer[1200] = 8'h78;
 buffer[1201] = 8'hcc;
 buffer[1202] = 8'h00;
 buffer[1203] = 8'hcc;
 buffer[1204] = 8'hcc;
 buffer[1205] = 8'hcc;
 buffer[1206] = 8'h7e;
 buffer[1207] = 8'h00;
 buffer[1208] = 8'h00;
 buffer[1209] = 8'he0;
 buffer[1210] = 8'h00;
 buffer[1211] = 8'hcc;
 buffer[1212] = 8'hcc;
 buffer[1213] = 8'hcc;
 buffer[1214] = 8'h7e;
 buffer[1215] = 8'h00;
 buffer[1216] = 8'h00;
 buffer[1217] = 8'hcc;
 buffer[1218] = 8'h00;
 buffer[1219] = 8'hcc;
 buffer[1220] = 8'hcc;
 buffer[1221] = 8'h7c;
 buffer[1222] = 8'h0c;
 buffer[1223] = 8'hf8;
 buffer[1224] = 8'hc3;
 buffer[1225] = 8'h18;
 buffer[1226] = 8'h3c;
 buffer[1227] = 8'h66;
 buffer[1228] = 8'h66;
 buffer[1229] = 8'h3c;
 buffer[1230] = 8'h18;
 buffer[1231] = 8'h00;
 buffer[1232] = 8'hcc;
 buffer[1233] = 8'h00;
 buffer[1234] = 8'hcc;
 buffer[1235] = 8'hcc;
 buffer[1236] = 8'hcc;
 buffer[1237] = 8'hcc;
 buffer[1238] = 8'h78;
 buffer[1239] = 8'h00;
 buffer[1240] = 8'h18;
 buffer[1241] = 8'h18;
 buffer[1242] = 8'h7e;
 buffer[1243] = 8'hc0;
 buffer[1244] = 8'hc0;
 buffer[1245] = 8'h7e;
 buffer[1246] = 8'h18;
 buffer[1247] = 8'h18;
 buffer[1248] = 8'h38;
 buffer[1249] = 8'h6c;
 buffer[1250] = 8'h64;
 buffer[1251] = 8'hf0;
 buffer[1252] = 8'h60;
 buffer[1253] = 8'he6;
 buffer[1254] = 8'hfc;
 buffer[1255] = 8'h00;
 buffer[1256] = 8'hcc;
 buffer[1257] = 8'hcc;
 buffer[1258] = 8'h78;
 buffer[1259] = 8'hfc;
 buffer[1260] = 8'h30;
 buffer[1261] = 8'hfc;
 buffer[1262] = 8'h30;
 buffer[1263] = 8'h30;
 buffer[1264] = 8'hf8;
 buffer[1265] = 8'hcc;
 buffer[1266] = 8'hcc;
 buffer[1267] = 8'hfa;
 buffer[1268] = 8'hc6;
 buffer[1269] = 8'hcf;
 buffer[1270] = 8'hc6;
 buffer[1271] = 8'hc7;
 buffer[1272] = 8'h0e;
 buffer[1273] = 8'h1b;
 buffer[1274] = 8'h18;
 buffer[1275] = 8'h3c;
 buffer[1276] = 8'h18;
 buffer[1277] = 8'h18;
 buffer[1278] = 8'hd8;
 buffer[1279] = 8'h70;
 buffer[1280] = 8'h1c;
 buffer[1281] = 8'h00;
 buffer[1282] = 8'h78;
 buffer[1283] = 8'h0c;
 buffer[1284] = 8'h7c;
 buffer[1285] = 8'hcc;
 buffer[1286] = 8'h7e;
 buffer[1287] = 8'h00;
 buffer[1288] = 8'h38;
 buffer[1289] = 8'h00;
 buffer[1290] = 8'h70;
 buffer[1291] = 8'h30;
 buffer[1292] = 8'h30;
 buffer[1293] = 8'h30;
 buffer[1294] = 8'h78;
 buffer[1295] = 8'h00;
 buffer[1296] = 8'h00;
 buffer[1297] = 8'h1c;
 buffer[1298] = 8'h00;
 buffer[1299] = 8'h78;
 buffer[1300] = 8'hcc;
 buffer[1301] = 8'hcc;
 buffer[1302] = 8'h78;
 buffer[1303] = 8'h00;
 buffer[1304] = 8'h00;
 buffer[1305] = 8'h1c;
 buffer[1306] = 8'h00;
 buffer[1307] = 8'hcc;
 buffer[1308] = 8'hcc;
 buffer[1309] = 8'hcc;
 buffer[1310] = 8'h7e;
 buffer[1311] = 8'h00;
 buffer[1312] = 8'h00;
 buffer[1313] = 8'hf8;
 buffer[1314] = 8'h00;
 buffer[1315] = 8'hf8;
 buffer[1316] = 8'hcc;
 buffer[1317] = 8'hcc;
 buffer[1318] = 8'hcc;
 buffer[1319] = 8'h00;
 buffer[1320] = 8'hfc;
 buffer[1321] = 8'h00;
 buffer[1322] = 8'hcc;
 buffer[1323] = 8'hec;
 buffer[1324] = 8'hfc;
 buffer[1325] = 8'hdc;
 buffer[1326] = 8'hcc;
 buffer[1327] = 8'h00;
 buffer[1328] = 8'h3c;
 buffer[1329] = 8'h6c;
 buffer[1330] = 8'h6c;
 buffer[1331] = 8'h3e;
 buffer[1332] = 8'h00;
 buffer[1333] = 8'h7e;
 buffer[1334] = 8'h00;
 buffer[1335] = 8'h00;
 buffer[1336] = 8'h38;
 buffer[1337] = 8'h6c;
 buffer[1338] = 8'h6c;
 buffer[1339] = 8'h38;
 buffer[1340] = 8'h00;
 buffer[1341] = 8'h7c;
 buffer[1342] = 8'h00;
 buffer[1343] = 8'h00;
 buffer[1344] = 8'h30;
 buffer[1345] = 8'h00;
 buffer[1346] = 8'h30;
 buffer[1347] = 8'h60;
 buffer[1348] = 8'hc0;
 buffer[1349] = 8'hcc;
 buffer[1350] = 8'h78;
 buffer[1351] = 8'h00;
 buffer[1352] = 8'h00;
 buffer[1353] = 8'h00;
 buffer[1354] = 8'h00;
 buffer[1355] = 8'hfc;
 buffer[1356] = 8'hc0;
 buffer[1357] = 8'hc0;
 buffer[1358] = 8'h00;
 buffer[1359] = 8'h00;
 buffer[1360] = 8'h00;
 buffer[1361] = 8'h00;
 buffer[1362] = 8'h00;
 buffer[1363] = 8'hfc;
 buffer[1364] = 8'h0c;
 buffer[1365] = 8'h0c;
 buffer[1366] = 8'h00;
 buffer[1367] = 8'h00;
 buffer[1368] = 8'hc3;
 buffer[1369] = 8'hc6;
 buffer[1370] = 8'hcc;
 buffer[1371] = 8'hde;
 buffer[1372] = 8'h33;
 buffer[1373] = 8'h66;
 buffer[1374] = 8'hcc;
 buffer[1375] = 8'h0f;
 buffer[1376] = 8'hc3;
 buffer[1377] = 8'hc6;
 buffer[1378] = 8'hcc;
 buffer[1379] = 8'hdb;
 buffer[1380] = 8'h37;
 buffer[1381] = 8'h6f;
 buffer[1382] = 8'hcf;
 buffer[1383] = 8'h03;
 buffer[1384] = 8'h18;
 buffer[1385] = 8'h18;
 buffer[1386] = 8'h00;
 buffer[1387] = 8'h18;
 buffer[1388] = 8'h18;
 buffer[1389] = 8'h18;
 buffer[1390] = 8'h18;
 buffer[1391] = 8'h00;
 buffer[1392] = 8'h00;
 buffer[1393] = 8'h33;
 buffer[1394] = 8'h66;
 buffer[1395] = 8'hcc;
 buffer[1396] = 8'h66;
 buffer[1397] = 8'h33;
 buffer[1398] = 8'h00;
 buffer[1399] = 8'h00;
 buffer[1400] = 8'h00;
 buffer[1401] = 8'hcc;
 buffer[1402] = 8'h66;
 buffer[1403] = 8'h33;
 buffer[1404] = 8'h66;
 buffer[1405] = 8'hcc;
 buffer[1406] = 8'h00;
 buffer[1407] = 8'h00;
 buffer[1408] = 8'h22;
 buffer[1409] = 8'h88;
 buffer[1410] = 8'h22;
 buffer[1411] = 8'h88;
 buffer[1412] = 8'h22;
 buffer[1413] = 8'h88;
 buffer[1414] = 8'h22;
 buffer[1415] = 8'h88;
 buffer[1416] = 8'h55;
 buffer[1417] = 8'haa;
 buffer[1418] = 8'h55;
 buffer[1419] = 8'haa;
 buffer[1420] = 8'h55;
 buffer[1421] = 8'haa;
 buffer[1422] = 8'h55;
 buffer[1423] = 8'haa;
 buffer[1424] = 8'hdb;
 buffer[1425] = 8'h77;
 buffer[1426] = 8'hdb;
 buffer[1427] = 8'hee;
 buffer[1428] = 8'hdb;
 buffer[1429] = 8'h77;
 buffer[1430] = 8'hdb;
 buffer[1431] = 8'hee;
 buffer[1432] = 8'h18;
 buffer[1433] = 8'h18;
 buffer[1434] = 8'h18;
 buffer[1435] = 8'h18;
 buffer[1436] = 8'h18;
 buffer[1437] = 8'h18;
 buffer[1438] = 8'h18;
 buffer[1439] = 8'h18;
 buffer[1440] = 8'h18;
 buffer[1441] = 8'h18;
 buffer[1442] = 8'h18;
 buffer[1443] = 8'h18;
 buffer[1444] = 8'hf8;
 buffer[1445] = 8'h18;
 buffer[1446] = 8'h18;
 buffer[1447] = 8'h18;
 buffer[1448] = 8'h18;
 buffer[1449] = 8'h18;
 buffer[1450] = 8'hf8;
 buffer[1451] = 8'h18;
 buffer[1452] = 8'hf8;
 buffer[1453] = 8'h18;
 buffer[1454] = 8'h18;
 buffer[1455] = 8'h18;
 buffer[1456] = 8'h36;
 buffer[1457] = 8'h36;
 buffer[1458] = 8'h36;
 buffer[1459] = 8'h36;
 buffer[1460] = 8'hf6;
 buffer[1461] = 8'h36;
 buffer[1462] = 8'h36;
 buffer[1463] = 8'h36;
 buffer[1464] = 8'h00;
 buffer[1465] = 8'h00;
 buffer[1466] = 8'h00;
 buffer[1467] = 8'h00;
 buffer[1468] = 8'hfe;
 buffer[1469] = 8'h36;
 buffer[1470] = 8'h36;
 buffer[1471] = 8'h36;
 buffer[1472] = 8'h00;
 buffer[1473] = 8'h00;
 buffer[1474] = 8'hf8;
 buffer[1475] = 8'h18;
 buffer[1476] = 8'hf8;
 buffer[1477] = 8'h18;
 buffer[1478] = 8'h18;
 buffer[1479] = 8'h18;
 buffer[1480] = 8'h36;
 buffer[1481] = 8'h36;
 buffer[1482] = 8'hf6;
 buffer[1483] = 8'h06;
 buffer[1484] = 8'hf6;
 buffer[1485] = 8'h36;
 buffer[1486] = 8'h36;
 buffer[1487] = 8'h36;
 buffer[1488] = 8'h36;
 buffer[1489] = 8'h36;
 buffer[1490] = 8'h36;
 buffer[1491] = 8'h36;
 buffer[1492] = 8'h36;
 buffer[1493] = 8'h36;
 buffer[1494] = 8'h36;
 buffer[1495] = 8'h36;
 buffer[1496] = 8'h00;
 buffer[1497] = 8'h00;
 buffer[1498] = 8'hfe;
 buffer[1499] = 8'h06;
 buffer[1500] = 8'hf6;
 buffer[1501] = 8'h36;
 buffer[1502] = 8'h36;
 buffer[1503] = 8'h36;
 buffer[1504] = 8'h36;
 buffer[1505] = 8'h36;
 buffer[1506] = 8'hf6;
 buffer[1507] = 8'h06;
 buffer[1508] = 8'hfe;
 buffer[1509] = 8'h00;
 buffer[1510] = 8'h00;
 buffer[1511] = 8'h00;
 buffer[1512] = 8'h36;
 buffer[1513] = 8'h36;
 buffer[1514] = 8'h36;
 buffer[1515] = 8'h36;
 buffer[1516] = 8'hfe;
 buffer[1517] = 8'h00;
 buffer[1518] = 8'h00;
 buffer[1519] = 8'h00;
 buffer[1520] = 8'h18;
 buffer[1521] = 8'h18;
 buffer[1522] = 8'hf8;
 buffer[1523] = 8'h18;
 buffer[1524] = 8'hf8;
 buffer[1525] = 8'h00;
 buffer[1526] = 8'h00;
 buffer[1527] = 8'h00;
 buffer[1528] = 8'h00;
 buffer[1529] = 8'h00;
 buffer[1530] = 8'h00;
 buffer[1531] = 8'h00;
 buffer[1532] = 8'hf8;
 buffer[1533] = 8'h18;
 buffer[1534] = 8'h18;
 buffer[1535] = 8'h18;
 buffer[1536] = 8'h18;
 buffer[1537] = 8'h18;
 buffer[1538] = 8'h18;
 buffer[1539] = 8'h18;
 buffer[1540] = 8'h1f;
 buffer[1541] = 8'h00;
 buffer[1542] = 8'h00;
 buffer[1543] = 8'h00;
 buffer[1544] = 8'h18;
 buffer[1545] = 8'h18;
 buffer[1546] = 8'h18;
 buffer[1547] = 8'h18;
 buffer[1548] = 8'hff;
 buffer[1549] = 8'h00;
 buffer[1550] = 8'h00;
 buffer[1551] = 8'h00;
 buffer[1552] = 8'h00;
 buffer[1553] = 8'h00;
 buffer[1554] = 8'h00;
 buffer[1555] = 8'h00;
 buffer[1556] = 8'hff;
 buffer[1557] = 8'h18;
 buffer[1558] = 8'h18;
 buffer[1559] = 8'h18;
 buffer[1560] = 8'h18;
 buffer[1561] = 8'h18;
 buffer[1562] = 8'h18;
 buffer[1563] = 8'h18;
 buffer[1564] = 8'h1f;
 buffer[1565] = 8'h18;
 buffer[1566] = 8'h18;
 buffer[1567] = 8'h18;
 buffer[1568] = 8'h00;
 buffer[1569] = 8'h00;
 buffer[1570] = 8'h00;
 buffer[1571] = 8'h00;
 buffer[1572] = 8'hff;
 buffer[1573] = 8'h00;
 buffer[1574] = 8'h00;
 buffer[1575] = 8'h00;
 buffer[1576] = 8'h18;
 buffer[1577] = 8'h18;
 buffer[1578] = 8'h18;
 buffer[1579] = 8'h18;
 buffer[1580] = 8'hff;
 buffer[1581] = 8'h18;
 buffer[1582] = 8'h18;
 buffer[1583] = 8'h18;
 buffer[1584] = 8'h18;
 buffer[1585] = 8'h18;
 buffer[1586] = 8'h1f;
 buffer[1587] = 8'h18;
 buffer[1588] = 8'h1f;
 buffer[1589] = 8'h18;
 buffer[1590] = 8'h18;
 buffer[1591] = 8'h18;
 buffer[1592] = 8'h36;
 buffer[1593] = 8'h36;
 buffer[1594] = 8'h36;
 buffer[1595] = 8'h36;
 buffer[1596] = 8'h37;
 buffer[1597] = 8'h36;
 buffer[1598] = 8'h36;
 buffer[1599] = 8'h36;
 buffer[1600] = 8'h36;
 buffer[1601] = 8'h36;
 buffer[1602] = 8'h37;
 buffer[1603] = 8'h30;
 buffer[1604] = 8'h3f;
 buffer[1605] = 8'h00;
 buffer[1606] = 8'h00;
 buffer[1607] = 8'h00;
 buffer[1608] = 8'h00;
 buffer[1609] = 8'h00;
 buffer[1610] = 8'h3f;
 buffer[1611] = 8'h30;
 buffer[1612] = 8'h37;
 buffer[1613] = 8'h36;
 buffer[1614] = 8'h36;
 buffer[1615] = 8'h36;
 buffer[1616] = 8'h36;
 buffer[1617] = 8'h36;
 buffer[1618] = 8'hf7;
 buffer[1619] = 8'h00;
 buffer[1620] = 8'hff;
 buffer[1621] = 8'h00;
 buffer[1622] = 8'h00;
 buffer[1623] = 8'h00;
 buffer[1624] = 8'h00;
 buffer[1625] = 8'h00;
 buffer[1626] = 8'hff;
 buffer[1627] = 8'h00;
 buffer[1628] = 8'hf7;
 buffer[1629] = 8'h36;
 buffer[1630] = 8'h36;
 buffer[1631] = 8'h36;
 buffer[1632] = 8'h36;
 buffer[1633] = 8'h36;
 buffer[1634] = 8'h37;
 buffer[1635] = 8'h30;
 buffer[1636] = 8'h37;
 buffer[1637] = 8'h36;
 buffer[1638] = 8'h36;
 buffer[1639] = 8'h36;
 buffer[1640] = 8'h00;
 buffer[1641] = 8'h00;
 buffer[1642] = 8'hff;
 buffer[1643] = 8'h00;
 buffer[1644] = 8'hff;
 buffer[1645] = 8'h00;
 buffer[1646] = 8'h00;
 buffer[1647] = 8'h00;
 buffer[1648] = 8'h36;
 buffer[1649] = 8'h36;
 buffer[1650] = 8'hf7;
 buffer[1651] = 8'h00;
 buffer[1652] = 8'hf7;
 buffer[1653] = 8'h36;
 buffer[1654] = 8'h36;
 buffer[1655] = 8'h36;
 buffer[1656] = 8'h18;
 buffer[1657] = 8'h18;
 buffer[1658] = 8'hff;
 buffer[1659] = 8'h00;
 buffer[1660] = 8'hff;
 buffer[1661] = 8'h00;
 buffer[1662] = 8'h00;
 buffer[1663] = 8'h00;
 buffer[1664] = 8'h36;
 buffer[1665] = 8'h36;
 buffer[1666] = 8'h36;
 buffer[1667] = 8'h36;
 buffer[1668] = 8'hff;
 buffer[1669] = 8'h00;
 buffer[1670] = 8'h00;
 buffer[1671] = 8'h00;
 buffer[1672] = 8'h00;
 buffer[1673] = 8'h00;
 buffer[1674] = 8'hff;
 buffer[1675] = 8'h00;
 buffer[1676] = 8'hff;
 buffer[1677] = 8'h18;
 buffer[1678] = 8'h18;
 buffer[1679] = 8'h18;
 buffer[1680] = 8'h00;
 buffer[1681] = 8'h00;
 buffer[1682] = 8'h00;
 buffer[1683] = 8'h00;
 buffer[1684] = 8'hff;
 buffer[1685] = 8'h36;
 buffer[1686] = 8'h36;
 buffer[1687] = 8'h36;
 buffer[1688] = 8'h36;
 buffer[1689] = 8'h36;
 buffer[1690] = 8'h36;
 buffer[1691] = 8'h36;
 buffer[1692] = 8'h3f;
 buffer[1693] = 8'h00;
 buffer[1694] = 8'h00;
 buffer[1695] = 8'h00;
 buffer[1696] = 8'h18;
 buffer[1697] = 8'h18;
 buffer[1698] = 8'h1f;
 buffer[1699] = 8'h18;
 buffer[1700] = 8'h1f;
 buffer[1701] = 8'h00;
 buffer[1702] = 8'h00;
 buffer[1703] = 8'h00;
 buffer[1704] = 8'h00;
 buffer[1705] = 8'h00;
 buffer[1706] = 8'h1f;
 buffer[1707] = 8'h18;
 buffer[1708] = 8'h1f;
 buffer[1709] = 8'h18;
 buffer[1710] = 8'h18;
 buffer[1711] = 8'h18;
 buffer[1712] = 8'h00;
 buffer[1713] = 8'h00;
 buffer[1714] = 8'h00;
 buffer[1715] = 8'h00;
 buffer[1716] = 8'h3f;
 buffer[1717] = 8'h36;
 buffer[1718] = 8'h36;
 buffer[1719] = 8'h36;
 buffer[1720] = 8'h36;
 buffer[1721] = 8'h36;
 buffer[1722] = 8'h36;
 buffer[1723] = 8'h36;
 buffer[1724] = 8'hff;
 buffer[1725] = 8'h36;
 buffer[1726] = 8'h36;
 buffer[1727] = 8'h36;
 buffer[1728] = 8'h18;
 buffer[1729] = 8'h18;
 buffer[1730] = 8'hff;
 buffer[1731] = 8'h18;
 buffer[1732] = 8'hff;
 buffer[1733] = 8'h18;
 buffer[1734] = 8'h18;
 buffer[1735] = 8'h18;
 buffer[1736] = 8'h18;
 buffer[1737] = 8'h18;
 buffer[1738] = 8'h18;
 buffer[1739] = 8'h18;
 buffer[1740] = 8'hf8;
 buffer[1741] = 8'h00;
 buffer[1742] = 8'h00;
 buffer[1743] = 8'h00;
 buffer[1744] = 8'h00;
 buffer[1745] = 8'h00;
 buffer[1746] = 8'h00;
 buffer[1747] = 8'h00;
 buffer[1748] = 8'h1f;
 buffer[1749] = 8'h18;
 buffer[1750] = 8'h18;
 buffer[1751] = 8'h18;
 buffer[1752] = 8'hff;
 buffer[1753] = 8'hff;
 buffer[1754] = 8'hff;
 buffer[1755] = 8'hff;
 buffer[1756] = 8'hff;
 buffer[1757] = 8'hff;
 buffer[1758] = 8'hff;
 buffer[1759] = 8'hff;
 buffer[1760] = 8'h00;
 buffer[1761] = 8'h00;
 buffer[1762] = 8'h00;
 buffer[1763] = 8'h00;
 buffer[1764] = 8'hff;
 buffer[1765] = 8'hff;
 buffer[1766] = 8'hff;
 buffer[1767] = 8'hff;
 buffer[1768] = 8'hf0;
 buffer[1769] = 8'hf0;
 buffer[1770] = 8'hf0;
 buffer[1771] = 8'hf0;
 buffer[1772] = 8'hf0;
 buffer[1773] = 8'hf0;
 buffer[1774] = 8'hf0;
 buffer[1775] = 8'hf0;
 buffer[1776] = 8'h0f;
 buffer[1777] = 8'h0f;
 buffer[1778] = 8'h0f;
 buffer[1779] = 8'h0f;
 buffer[1780] = 8'h0f;
 buffer[1781] = 8'h0f;
 buffer[1782] = 8'h0f;
 buffer[1783] = 8'h0f;
 buffer[1784] = 8'hff;
 buffer[1785] = 8'hff;
 buffer[1786] = 8'hff;
 buffer[1787] = 8'hff;
 buffer[1788] = 8'h00;
 buffer[1789] = 8'h00;
 buffer[1790] = 8'h00;
 buffer[1791] = 8'h00;
 buffer[1792] = 8'h00;
 buffer[1793] = 8'h00;
 buffer[1794] = 8'h76;
 buffer[1795] = 8'hdc;
 buffer[1796] = 8'hc8;
 buffer[1797] = 8'hdc;
 buffer[1798] = 8'h76;
 buffer[1799] = 8'h00;
 buffer[1800] = 8'h00;
 buffer[1801] = 8'h78;
 buffer[1802] = 8'hcc;
 buffer[1803] = 8'hf8;
 buffer[1804] = 8'hcc;
 buffer[1805] = 8'hf8;
 buffer[1806] = 8'hc0;
 buffer[1807] = 8'hc0;
 buffer[1808] = 8'h00;
 buffer[1809] = 8'hfc;
 buffer[1810] = 8'hcc;
 buffer[1811] = 8'hc0;
 buffer[1812] = 8'hc0;
 buffer[1813] = 8'hc0;
 buffer[1814] = 8'hc0;
 buffer[1815] = 8'h00;
 buffer[1816] = 8'h00;
 buffer[1817] = 8'hfe;
 buffer[1818] = 8'h6c;
 buffer[1819] = 8'h6c;
 buffer[1820] = 8'h6c;
 buffer[1821] = 8'h6c;
 buffer[1822] = 8'h6c;
 buffer[1823] = 8'h00;
 buffer[1824] = 8'hfc;
 buffer[1825] = 8'hcc;
 buffer[1826] = 8'h60;
 buffer[1827] = 8'h30;
 buffer[1828] = 8'h60;
 buffer[1829] = 8'hcc;
 buffer[1830] = 8'hfc;
 buffer[1831] = 8'h00;
 buffer[1832] = 8'h00;
 buffer[1833] = 8'h00;
 buffer[1834] = 8'h7e;
 buffer[1835] = 8'hd8;
 buffer[1836] = 8'hd8;
 buffer[1837] = 8'hd8;
 buffer[1838] = 8'h70;
 buffer[1839] = 8'h00;
 buffer[1840] = 8'h00;
 buffer[1841] = 8'h66;
 buffer[1842] = 8'h66;
 buffer[1843] = 8'h66;
 buffer[1844] = 8'h66;
 buffer[1845] = 8'h7c;
 buffer[1846] = 8'h60;
 buffer[1847] = 8'hc0;
 buffer[1848] = 8'h00;
 buffer[1849] = 8'h76;
 buffer[1850] = 8'hdc;
 buffer[1851] = 8'h18;
 buffer[1852] = 8'h18;
 buffer[1853] = 8'h18;
 buffer[1854] = 8'h18;
 buffer[1855] = 8'h00;
 buffer[1856] = 8'hfc;
 buffer[1857] = 8'h30;
 buffer[1858] = 8'h78;
 buffer[1859] = 8'hcc;
 buffer[1860] = 8'hcc;
 buffer[1861] = 8'h78;
 buffer[1862] = 8'h30;
 buffer[1863] = 8'hfc;
 buffer[1864] = 8'h38;
 buffer[1865] = 8'h6c;
 buffer[1866] = 8'hc6;
 buffer[1867] = 8'hfe;
 buffer[1868] = 8'hc6;
 buffer[1869] = 8'h6c;
 buffer[1870] = 8'h38;
 buffer[1871] = 8'h00;
 buffer[1872] = 8'h38;
 buffer[1873] = 8'h6c;
 buffer[1874] = 8'hc6;
 buffer[1875] = 8'hc6;
 buffer[1876] = 8'h6c;
 buffer[1877] = 8'h6c;
 buffer[1878] = 8'hee;
 buffer[1879] = 8'h00;
 buffer[1880] = 8'h1c;
 buffer[1881] = 8'h30;
 buffer[1882] = 8'h18;
 buffer[1883] = 8'h7c;
 buffer[1884] = 8'hcc;
 buffer[1885] = 8'hcc;
 buffer[1886] = 8'h78;
 buffer[1887] = 8'h00;
 buffer[1888] = 8'h00;
 buffer[1889] = 8'h00;
 buffer[1890] = 8'h7e;
 buffer[1891] = 8'hdb;
 buffer[1892] = 8'hdb;
 buffer[1893] = 8'h7e;
 buffer[1894] = 8'h00;
 buffer[1895] = 8'h00;
 buffer[1896] = 8'h06;
 buffer[1897] = 8'h0c;
 buffer[1898] = 8'h7e;
 buffer[1899] = 8'hdb;
 buffer[1900] = 8'hdb;
 buffer[1901] = 8'h7e;
 buffer[1902] = 8'h60;
 buffer[1903] = 8'hc0;
 buffer[1904] = 8'h38;
 buffer[1905] = 8'h60;
 buffer[1906] = 8'hc0;
 buffer[1907] = 8'hf8;
 buffer[1908] = 8'hc0;
 buffer[1909] = 8'h60;
 buffer[1910] = 8'h38;
 buffer[1911] = 8'h00;
 buffer[1912] = 8'h78;
 buffer[1913] = 8'hcc;
 buffer[1914] = 8'hcc;
 buffer[1915] = 8'hcc;
 buffer[1916] = 8'hcc;
 buffer[1917] = 8'hcc;
 buffer[1918] = 8'hcc;
 buffer[1919] = 8'h00;
 buffer[1920] = 8'h00;
 buffer[1921] = 8'hfc;
 buffer[1922] = 8'h00;
 buffer[1923] = 8'hfc;
 buffer[1924] = 8'h00;
 buffer[1925] = 8'hfc;
 buffer[1926] = 8'h00;
 buffer[1927] = 8'h00;
 buffer[1928] = 8'h30;
 buffer[1929] = 8'h30;
 buffer[1930] = 8'hfc;
 buffer[1931] = 8'h30;
 buffer[1932] = 8'h30;
 buffer[1933] = 8'h00;
 buffer[1934] = 8'hfc;
 buffer[1935] = 8'h00;
 buffer[1936] = 8'h60;
 buffer[1937] = 8'h30;
 buffer[1938] = 8'h18;
 buffer[1939] = 8'h30;
 buffer[1940] = 8'h60;
 buffer[1941] = 8'h00;
 buffer[1942] = 8'hfc;
 buffer[1943] = 8'h00;
 buffer[1944] = 8'h18;
 buffer[1945] = 8'h30;
 buffer[1946] = 8'h60;
 buffer[1947] = 8'h30;
 buffer[1948] = 8'h18;
 buffer[1949] = 8'h00;
 buffer[1950] = 8'hfc;
 buffer[1951] = 8'h00;
 buffer[1952] = 8'h0e;
 buffer[1953] = 8'h1b;
 buffer[1954] = 8'h1b;
 buffer[1955] = 8'h18;
 buffer[1956] = 8'h18;
 buffer[1957] = 8'h18;
 buffer[1958] = 8'h18;
 buffer[1959] = 8'h18;
 buffer[1960] = 8'h18;
 buffer[1961] = 8'h18;
 buffer[1962] = 8'h18;
 buffer[1963] = 8'h18;
 buffer[1964] = 8'h18;
 buffer[1965] = 8'hd8;
 buffer[1966] = 8'hd8;
 buffer[1967] = 8'h70;
 buffer[1968] = 8'h30;
 buffer[1969] = 8'h30;
 buffer[1970] = 8'h00;
 buffer[1971] = 8'hfc;
 buffer[1972] = 8'h00;
 buffer[1973] = 8'h30;
 buffer[1974] = 8'h30;
 buffer[1975] = 8'h00;
 buffer[1976] = 8'h00;
 buffer[1977] = 8'h76;
 buffer[1978] = 8'hdc;
 buffer[1979] = 8'h00;
 buffer[1980] = 8'h76;
 buffer[1981] = 8'hdc;
 buffer[1982] = 8'h00;
 buffer[1983] = 8'h00;
 buffer[1984] = 8'h38;
 buffer[1985] = 8'h6c;
 buffer[1986] = 8'h6c;
 buffer[1987] = 8'h38;
 buffer[1988] = 8'h00;
 buffer[1989] = 8'h00;
 buffer[1990] = 8'h00;
 buffer[1991] = 8'h00;
 buffer[1992] = 8'h00;
 buffer[1993] = 8'h00;
 buffer[1994] = 8'h00;
 buffer[1995] = 8'h18;
 buffer[1996] = 8'h18;
 buffer[1997] = 8'h00;
 buffer[1998] = 8'h00;
 buffer[1999] = 8'h00;
 buffer[2000] = 8'h00;
 buffer[2001] = 8'h00;
 buffer[2002] = 8'h00;
 buffer[2003] = 8'h00;
 buffer[2004] = 8'h18;
 buffer[2005] = 8'h00;
 buffer[2006] = 8'h00;
 buffer[2007] = 8'h00;
 buffer[2008] = 8'h0f;
 buffer[2009] = 8'h0c;
 buffer[2010] = 8'h0c;
 buffer[2011] = 8'h0c;
 buffer[2012] = 8'hec;
 buffer[2013] = 8'h6c;
 buffer[2014] = 8'h3c;
 buffer[2015] = 8'h1c;
 buffer[2016] = 8'h78;
 buffer[2017] = 8'h6c;
 buffer[2018] = 8'h6c;
 buffer[2019] = 8'h6c;
 buffer[2020] = 8'h6c;
 buffer[2021] = 8'h00;
 buffer[2022] = 8'h00;
 buffer[2023] = 8'h00;
 buffer[2024] = 8'h70;
 buffer[2025] = 8'h18;
 buffer[2026] = 8'h30;
 buffer[2027] = 8'h60;
 buffer[2028] = 8'h78;
 buffer[2029] = 8'h00;
 buffer[2030] = 8'h00;
 buffer[2031] = 8'h00;
 buffer[2032] = 8'h00;
 buffer[2033] = 8'h00;
 buffer[2034] = 8'h3c;
 buffer[2035] = 8'h3c;
 buffer[2036] = 8'h3c;
 buffer[2037] = 8'h3c;
 buffer[2038] = 8'h00;
 buffer[2039] = 8'h00;
 buffer[2040] = 8'h00;
 buffer[2041] = 8'h00;
 buffer[2042] = 8'h00;
 buffer[2043] = 8'h00;
 buffer[2044] = 8'h00;
 buffer[2045] = 8'h00;
 buffer[2046] = 8'h00;
 buffer[2047] = 8'h00;
end

endmodule

module M_terminal_mem_terminal(
input      [9:0]                in_terminal_addr0,
output reg  [7:0]     out_terminal_rdata0,
output reg  [7:0]     out_terminal_rdata1,
input      [0:0]             in_terminal_wenable1,
input      [7:0]                 in_terminal_wdata1,
input      [9:0]                in_terminal_addr1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[639:0];
always @(posedge clock0) begin
  out_terminal_rdata0 <= buffer[in_terminal_addr0];
end
always @(posedge clock1) begin
  if (in_terminal_wenable1) begin
    buffer[in_terminal_addr1] <= in_terminal_wdata1;
  end
end

endmodule

module M_terminal_mem_terminal_copy(
input      [9:0]                in_terminal_copy_addr0,
output reg  [7:0]     out_terminal_copy_rdata0,
output reg  [7:0]     out_terminal_copy_rdata1,
input      [0:0]             in_terminal_copy_wenable1,
input      [7:0]                 in_terminal_copy_wdata1,
input      [9:0]                in_terminal_copy_addr1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[639:0];
always @(posedge clock0) begin
  out_terminal_copy_rdata0 <= buffer[in_terminal_copy_addr0];
end
always @(posedge clock1) begin
  if (in_terminal_copy_wenable1) begin
    buffer[in_terminal_copy_addr1] <= in_terminal_copy_wdata1;
  end
end

endmodule

module M_terminal (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_terminal_character,
in_terminal_write,
in_showterminal,
in_timer1hz,
out_pix_red,
out_pix_green,
out_pix_blue,
out_terminal_display,
out_terminal_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [7:0] in_terminal_character;
input  [1:0] in_terminal_write;
input  [0:0] in_showterminal;
input  [0:0] in_timer1hz;
output  [1:0] out_pix_red;
output  [1:0] out_pix_green;
output  [1:0] out_pix_blue;
output  [0:0] out_terminal_display;
output  [1:0] out_terminal_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [7:0] _w_mem_characterGenerator8x8_rdata;
wire  [7:0] _w_mem_terminal_rdata0;
wire  [7:0] _w_mem_terminal_copy_rdata0;
reg  [9:0] _t_terminal_addr0;
reg  [0:0] _t_terminal_wenable1;
reg  [7:0] _t_terminal_wdata1;
reg  [9:0] _t_terminal_addr1;
reg  [9:0] _t_terminal_copy_addr0;
reg  [0:0] _t_terminal_copy_wenable1;
reg  [7:0] _t_terminal_copy_wdata1;
reg  [9:0] _t_terminal_copy_addr1;
wire  [6:0] _w_xterminalpos;
wire  [9:0] _w_yterminalpos;
wire  [0:0] _w_is_cursor;
wire  [2:0] _w_xinterminal;
wire  [2:0] _w_yinterminal;
wire  [0:0] _w_terminalpixel;

reg  [10:0] _d_characterGenerator8x8_addr;
reg  [10:0] _q_characterGenerator8x8_addr;
reg  [6:0] _d_terminal_x;
reg  [6:0] _q_terminal_x;
reg  [2:0] _d_terminal_y;
reg  [2:0] _q_terminal_y;
reg  [9:0] _d_terminal_scroll;
reg  [9:0] _q_terminal_scroll;
reg  [1:0] _d_pix_red,_q_pix_red;
reg  [1:0] _d_pix_green,_q_pix_green;
reg  [1:0] _d_pix_blue,_q_pix_blue;
reg  [0:0] _d_terminal_display,_q_terminal_display;
reg  [1:0] _d_terminal_active,_q_terminal_active;
reg  [3:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_terminal_display = _d_terminal_display;
assign out_terminal_active = _q_terminal_active;
assign out_done = (_q_index == 11);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_characterGenerator8x8_addr <= 0;
_q_terminal_x <= 0;
_q_terminal_y <= 7;
_q_terminal_scroll <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_characterGenerator8x8_addr <= _d_characterGenerator8x8_addr;
_q_terminal_x <= _d_terminal_x;
_q_terminal_y <= _d_terminal_y;
_q_terminal_scroll <= _d_terminal_scroll;
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_terminal_display <= _d_terminal_display;
_q_terminal_active <= _d_terminal_active;
_q_index <= _d_index;
  end
end


M_terminal_mem_characterGenerator8x8 __mem__characterGenerator8x8(
.clock(clock),
.in_characterGenerator8x8_addr(_d_characterGenerator8x8_addr),
.out_characterGenerator8x8_rdata(_w_mem_characterGenerator8x8_rdata)
);
M_terminal_mem_terminal __mem__terminal(
.clock0(clock),
.clock1(clock),
.in_terminal_addr0(_t_terminal_addr0),
.in_terminal_wenable1(_t_terminal_wenable1),
.in_terminal_wdata1(_t_terminal_wdata1),
.in_terminal_addr1(_t_terminal_addr1),
.out_terminal_rdata0(_w_mem_terminal_rdata0)
);
M_terminal_mem_terminal_copy __mem__terminal_copy(
.clock0(clock),
.clock1(clock),
.in_terminal_copy_addr0(_t_terminal_copy_addr0),
.in_terminal_copy_wenable1(_t_terminal_copy_wenable1),
.in_terminal_copy_wdata1(_t_terminal_copy_wdata1),
.in_terminal_copy_addr1(_t_terminal_copy_addr1),
.out_terminal_copy_rdata0(_w_mem_terminal_copy_rdata0)
);

assign _w_terminalpixel = _w_mem_characterGenerator8x8_rdata[7-_w_xinterminal+:1];
assign _w_yinterminal = (in_pix_y)&7;
assign _w_xinterminal = (in_pix_x)&7;
assign _w_is_cursor = (_w_xterminalpos==_d_terminal_x)&&(((in_pix_y-416)>>3)==_d_terminal_y);
assign _w_yterminalpos = ((in_pix_vblank?0:in_pix_y-416)>>3)*80;
assign _w_xterminalpos = (in_pix_active?in_pix_x+2:0)>>3;

always @* begin
_d_characterGenerator8x8_addr = _q_characterGenerator8x8_addr;
_d_terminal_x = _q_terminal_x;
_d_terminal_y = _q_terminal_y;
_d_terminal_scroll = _q_terminal_scroll;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_terminal_display = _q_terminal_display;
_d_terminal_active = _q_terminal_active;
_d_index = _q_index;
_t_terminal_addr0 = 0;
_t_terminal_wenable1 = 0;
_t_terminal_wdata1 = 0;
_t_terminal_addr1 = 0;
_t_terminal_copy_addr0 = 0;
_t_terminal_copy_wenable1 = 0;
_t_terminal_copy_wdata1 = 0;
_t_terminal_copy_addr1 = 0;
// _always_pre
_t_terminal_addr0 = _w_xterminalpos+_w_yterminalpos;
_t_terminal_wenable1 = 1;
_t_terminal_copy_wenable1 = 1;
_d_characterGenerator8x8_addr = _w_mem_terminal_rdata0*8+_w_yinterminal;
_d_terminal_display = in_pix_active&&in_showterminal&&(in_pix_y>415);
_d_pix_red = (_w_terminalpixel)?((_w_is_cursor&&in_timer1hz)?0:3):((_w_is_cursor&&in_timer1hz)?3:0);
_d_pix_green = (_w_terminalpixel)?((_w_is_cursor&&in_timer1hz)?0:3):((_w_is_cursor&&in_timer1hz)?3:0);
_d_pix_blue = 3;
_d_index = 11;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_characterGenerator8x8_addr = 0;
_t_terminal_addr0 = 0;
_t_terminal_wenable1 = 0;
_t_terminal_wdata1 = 0;
_t_terminal_addr1 = 0;
_t_terminal_copy_addr0 = 0;
_t_terminal_copy_wenable1 = 0;
_t_terminal_copy_wdata1 = 0;
_t_terminal_copy_addr1 = 0;
_d_terminal_x = 0;
_d_terminal_y = 7;
_d_terminal_scroll = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (_q_terminal_active)
  0: begin
// __block_6_case
// __block_7
  case (in_terminal_write)
  1: begin
// __block_9_case
// __block_10
  case (in_terminal_character)
  8: begin
// __block_12_case
// __block_13
if (_q_terminal_x!=0) begin
// __block_14
// __block_16
_d_terminal_x = _q_terminal_x-1;
_t_terminal_addr1 = _d_terminal_x+_q_terminal_y*80;
_t_terminal_wdata1 = 0;
_t_terminal_copy_addr1 = _d_terminal_x+_q_terminal_y*80;
_t_terminal_copy_wdata1 = 0;
// __block_17
end else begin
// __block_15
end
// __block_18
// __block_19
  end
  10: begin
// __block_20_case
// __block_21
_d_terminal_active = 1;
// __block_22
  end
  13: begin
// __block_23_case
// __block_24
_d_terminal_x = 0;
// __block_25
  end
  default: begin
// __block_26_case
// __block_27
_t_terminal_addr1 = _q_terminal_x+_q_terminal_y*80;
_t_terminal_wdata1 = in_terminal_character;
_t_terminal_copy_addr1 = _q_terminal_x+_q_terminal_y*80;
_t_terminal_copy_wdata1 = in_terminal_character;
_d_terminal_active = (_q_terminal_x==79)?1:0;
_d_terminal_x = (_q_terminal_x==79)?0:_q_terminal_x+1;
// __block_28
  end
endcase
// __block_11
// __block_29
  end
  2: begin
// __block_30_case
// __block_31
_d_terminal_active = 2;
// __block_32
  end
endcase
// __block_8
// __block_33
_d_index = 1;
  end
  1: begin
// __block_34_case
// __block_35
_d_terminal_scroll = 0;
_d_index = 3;
  end
  2: begin
// __block_49_case
// __block_50
_d_terminal_scroll = 0;
_d_index = 4;
  end
endcase
end else begin
_d_index = 2;
end
end
3: begin
// __block_36
_d_index = 5;
end
4: begin
// __block_51
_d_index = 6;
end
2: begin
// __block_3
_d_index = 11;
end
5: begin
// __while__block_37
if (_q_terminal_scroll<560) begin
// __block_38
// __block_40
_t_terminal_copy_addr0 = _q_terminal_scroll+80;
_d_index = 10;
end else begin
_d_index = 7;
end
end
6: begin
// __while__block_52
if (_q_terminal_scroll<640) begin
// __block_53
// __block_55
_t_terminal_addr1 = _q_terminal_scroll;
_t_terminal_wdata1 = 0;
_t_terminal_copy_addr1 = _q_terminal_scroll;
_t_terminal_copy_wdata1 = 0;
_d_terminal_scroll = _q_terminal_scroll+1;
// __block_56
_d_index = 6;
end else begin
_d_index = 8;
end
end
10: begin
// __block_41
_t_terminal_addr1 = _q_terminal_scroll;
_t_terminal_wdata1 = _w_mem_terminal_copy_rdata0;
_t_terminal_copy_addr1 = _q_terminal_scroll;
_t_terminal_copy_wdata1 = _w_mem_terminal_copy_rdata0;
_d_terminal_scroll = _q_terminal_scroll+1;
// __block_42
_d_index = 5;
end
7: begin
// __while__block_43
if (_q_terminal_scroll<640) begin
// __block_44
// __block_46
_t_terminal_addr1 = _q_terminal_scroll;
_t_terminal_wdata1 = 0;
_t_terminal_copy_addr1 = _q_terminal_scroll;
_t_terminal_copy_wdata1 = 0;
_d_terminal_scroll = _q_terminal_scroll+1;
// __block_47
_d_index = 7;
end else begin
_d_index = 9;
end
end
8: begin
// __block_54
_d_terminal_x = 0;
_d_terminal_y = 7;
_d_terminal_active = 0;
// __block_57
_d_index = 1;
end
9: begin
// __block_45
_d_terminal_active = 0;
// __block_48
_d_index = 1;
end
11: begin // end of terminal
end
default: begin 
_d_index = 11;
 end
endcase
end
endmodule


module M_character_map_mem_characterGenerator8x16(
input                  [11:0] in_characterGenerator8x16_addr,
output reg  [7:0] out_characterGenerator8x16_rdata,
input                                   clock
);
reg  [7:0] buffer[4095:0];
always @(posedge clock) begin
   out_characterGenerator8x16_rdata <= buffer[in_characterGenerator8x16_addr];
end
initial begin
 buffer[0] = 8'h00;
 buffer[1] = 8'h00;
 buffer[2] = 8'h00;
 buffer[3] = 8'h00;
 buffer[4] = 8'h00;
 buffer[5] = 8'h00;
 buffer[6] = 8'h00;
 buffer[7] = 8'h00;
 buffer[8] = 8'h00;
 buffer[9] = 8'h00;
 buffer[10] = 8'h00;
 buffer[11] = 8'h00;
 buffer[12] = 8'h00;
 buffer[13] = 8'h00;
 buffer[14] = 8'h00;
 buffer[15] = 8'h00;
 buffer[16] = 8'h00;
 buffer[17] = 8'h00;
 buffer[18] = 8'h7e;
 buffer[19] = 8'h81;
 buffer[20] = 8'ha5;
 buffer[21] = 8'h81;
 buffer[22] = 8'h81;
 buffer[23] = 8'hbd;
 buffer[24] = 8'h99;
 buffer[25] = 8'h81;
 buffer[26] = 8'h81;
 buffer[27] = 8'h7e;
 buffer[28] = 8'h00;
 buffer[29] = 8'h00;
 buffer[30] = 8'h00;
 buffer[31] = 8'h00;
 buffer[32] = 8'h00;
 buffer[33] = 8'h00;
 buffer[34] = 8'h7e;
 buffer[35] = 8'hff;
 buffer[36] = 8'hdb;
 buffer[37] = 8'hff;
 buffer[38] = 8'hff;
 buffer[39] = 8'hc3;
 buffer[40] = 8'he7;
 buffer[41] = 8'hff;
 buffer[42] = 8'hff;
 buffer[43] = 8'h7e;
 buffer[44] = 8'h00;
 buffer[45] = 8'h00;
 buffer[46] = 8'h00;
 buffer[47] = 8'h00;
 buffer[48] = 8'h00;
 buffer[49] = 8'h00;
 buffer[50] = 8'h00;
 buffer[51] = 8'h00;
 buffer[52] = 8'h6c;
 buffer[53] = 8'hfe;
 buffer[54] = 8'hfe;
 buffer[55] = 8'hfe;
 buffer[56] = 8'hfe;
 buffer[57] = 8'h7c;
 buffer[58] = 8'h38;
 buffer[59] = 8'h10;
 buffer[60] = 8'h00;
 buffer[61] = 8'h00;
 buffer[62] = 8'h00;
 buffer[63] = 8'h00;
 buffer[64] = 8'h00;
 buffer[65] = 8'h00;
 buffer[66] = 8'h00;
 buffer[67] = 8'h00;
 buffer[68] = 8'h10;
 buffer[69] = 8'h38;
 buffer[70] = 8'h7c;
 buffer[71] = 8'hfe;
 buffer[72] = 8'h7c;
 buffer[73] = 8'h38;
 buffer[74] = 8'h10;
 buffer[75] = 8'h00;
 buffer[76] = 8'h00;
 buffer[77] = 8'h00;
 buffer[78] = 8'h00;
 buffer[79] = 8'h00;
 buffer[80] = 8'h00;
 buffer[81] = 8'h00;
 buffer[82] = 8'h00;
 buffer[83] = 8'h18;
 buffer[84] = 8'h3c;
 buffer[85] = 8'h3c;
 buffer[86] = 8'he7;
 buffer[87] = 8'he7;
 buffer[88] = 8'he7;
 buffer[89] = 8'h18;
 buffer[90] = 8'h18;
 buffer[91] = 8'h3c;
 buffer[92] = 8'h00;
 buffer[93] = 8'h00;
 buffer[94] = 8'h00;
 buffer[95] = 8'h00;
 buffer[96] = 8'h00;
 buffer[97] = 8'h00;
 buffer[98] = 8'h00;
 buffer[99] = 8'h18;
 buffer[100] = 8'h3c;
 buffer[101] = 8'h7e;
 buffer[102] = 8'hff;
 buffer[103] = 8'hff;
 buffer[104] = 8'h7e;
 buffer[105] = 8'h18;
 buffer[106] = 8'h18;
 buffer[107] = 8'h3c;
 buffer[108] = 8'h00;
 buffer[109] = 8'h00;
 buffer[110] = 8'h00;
 buffer[111] = 8'h00;
 buffer[112] = 8'h00;
 buffer[113] = 8'h00;
 buffer[114] = 8'h00;
 buffer[115] = 8'h00;
 buffer[116] = 8'h00;
 buffer[117] = 8'h00;
 buffer[118] = 8'h18;
 buffer[119] = 8'h3c;
 buffer[120] = 8'h3c;
 buffer[121] = 8'h18;
 buffer[122] = 8'h00;
 buffer[123] = 8'h00;
 buffer[124] = 8'h00;
 buffer[125] = 8'h00;
 buffer[126] = 8'h00;
 buffer[127] = 8'h00;
 buffer[128] = 8'hff;
 buffer[129] = 8'hff;
 buffer[130] = 8'hff;
 buffer[131] = 8'hff;
 buffer[132] = 8'hff;
 buffer[133] = 8'hff;
 buffer[134] = 8'he7;
 buffer[135] = 8'hc3;
 buffer[136] = 8'hc3;
 buffer[137] = 8'he7;
 buffer[138] = 8'hff;
 buffer[139] = 8'hff;
 buffer[140] = 8'hff;
 buffer[141] = 8'hff;
 buffer[142] = 8'hff;
 buffer[143] = 8'hff;
 buffer[144] = 8'h00;
 buffer[145] = 8'h00;
 buffer[146] = 8'h00;
 buffer[147] = 8'h00;
 buffer[148] = 8'h00;
 buffer[149] = 8'h3c;
 buffer[150] = 8'h66;
 buffer[151] = 8'h42;
 buffer[152] = 8'h42;
 buffer[153] = 8'h66;
 buffer[154] = 8'h3c;
 buffer[155] = 8'h00;
 buffer[156] = 8'h00;
 buffer[157] = 8'h00;
 buffer[158] = 8'h00;
 buffer[159] = 8'h00;
 buffer[160] = 8'hff;
 buffer[161] = 8'hff;
 buffer[162] = 8'hff;
 buffer[163] = 8'hff;
 buffer[164] = 8'hff;
 buffer[165] = 8'hc3;
 buffer[166] = 8'h99;
 buffer[167] = 8'hbd;
 buffer[168] = 8'hbd;
 buffer[169] = 8'h99;
 buffer[170] = 8'hc3;
 buffer[171] = 8'hff;
 buffer[172] = 8'hff;
 buffer[173] = 8'hff;
 buffer[174] = 8'hff;
 buffer[175] = 8'hff;
 buffer[176] = 8'h00;
 buffer[177] = 8'h00;
 buffer[178] = 8'h1e;
 buffer[179] = 8'h0e;
 buffer[180] = 8'h1a;
 buffer[181] = 8'h32;
 buffer[182] = 8'h78;
 buffer[183] = 8'hcc;
 buffer[184] = 8'hcc;
 buffer[185] = 8'hcc;
 buffer[186] = 8'hcc;
 buffer[187] = 8'h78;
 buffer[188] = 8'h00;
 buffer[189] = 8'h00;
 buffer[190] = 8'h00;
 buffer[191] = 8'h00;
 buffer[192] = 8'h00;
 buffer[193] = 8'h00;
 buffer[194] = 8'h3c;
 buffer[195] = 8'h66;
 buffer[196] = 8'h66;
 buffer[197] = 8'h66;
 buffer[198] = 8'h66;
 buffer[199] = 8'h3c;
 buffer[200] = 8'h18;
 buffer[201] = 8'h7e;
 buffer[202] = 8'h18;
 buffer[203] = 8'h18;
 buffer[204] = 8'h00;
 buffer[205] = 8'h00;
 buffer[206] = 8'h00;
 buffer[207] = 8'h00;
 buffer[208] = 8'h00;
 buffer[209] = 8'h00;
 buffer[210] = 8'h3f;
 buffer[211] = 8'h33;
 buffer[212] = 8'h3f;
 buffer[213] = 8'h30;
 buffer[214] = 8'h30;
 buffer[215] = 8'h30;
 buffer[216] = 8'h30;
 buffer[217] = 8'h70;
 buffer[218] = 8'hf0;
 buffer[219] = 8'he0;
 buffer[220] = 8'h00;
 buffer[221] = 8'h00;
 buffer[222] = 8'h00;
 buffer[223] = 8'h00;
 buffer[224] = 8'h00;
 buffer[225] = 8'h00;
 buffer[226] = 8'h7f;
 buffer[227] = 8'h63;
 buffer[228] = 8'h7f;
 buffer[229] = 8'h63;
 buffer[230] = 8'h63;
 buffer[231] = 8'h63;
 buffer[232] = 8'h63;
 buffer[233] = 8'h67;
 buffer[234] = 8'he7;
 buffer[235] = 8'he6;
 buffer[236] = 8'hc0;
 buffer[237] = 8'h00;
 buffer[238] = 8'h00;
 buffer[239] = 8'h00;
 buffer[240] = 8'h00;
 buffer[241] = 8'h00;
 buffer[242] = 8'h00;
 buffer[243] = 8'h18;
 buffer[244] = 8'h18;
 buffer[245] = 8'hdb;
 buffer[246] = 8'h3c;
 buffer[247] = 8'he7;
 buffer[248] = 8'h3c;
 buffer[249] = 8'hdb;
 buffer[250] = 8'h18;
 buffer[251] = 8'h18;
 buffer[252] = 8'h00;
 buffer[253] = 8'h00;
 buffer[254] = 8'h00;
 buffer[255] = 8'h00;
 buffer[256] = 8'h00;
 buffer[257] = 8'h80;
 buffer[258] = 8'hc0;
 buffer[259] = 8'he0;
 buffer[260] = 8'hf0;
 buffer[261] = 8'hf8;
 buffer[262] = 8'hfe;
 buffer[263] = 8'hf8;
 buffer[264] = 8'hf0;
 buffer[265] = 8'he0;
 buffer[266] = 8'hc0;
 buffer[267] = 8'h80;
 buffer[268] = 8'h00;
 buffer[269] = 8'h00;
 buffer[270] = 8'h00;
 buffer[271] = 8'h00;
 buffer[272] = 8'h00;
 buffer[273] = 8'h02;
 buffer[274] = 8'h06;
 buffer[275] = 8'h0e;
 buffer[276] = 8'h1e;
 buffer[277] = 8'h3e;
 buffer[278] = 8'hfe;
 buffer[279] = 8'h3e;
 buffer[280] = 8'h1e;
 buffer[281] = 8'h0e;
 buffer[282] = 8'h06;
 buffer[283] = 8'h02;
 buffer[284] = 8'h00;
 buffer[285] = 8'h00;
 buffer[286] = 8'h00;
 buffer[287] = 8'h00;
 buffer[288] = 8'h00;
 buffer[289] = 8'h00;
 buffer[290] = 8'h18;
 buffer[291] = 8'h3c;
 buffer[292] = 8'h7e;
 buffer[293] = 8'h18;
 buffer[294] = 8'h18;
 buffer[295] = 8'h18;
 buffer[296] = 8'h7e;
 buffer[297] = 8'h3c;
 buffer[298] = 8'h18;
 buffer[299] = 8'h00;
 buffer[300] = 8'h00;
 buffer[301] = 8'h00;
 buffer[302] = 8'h00;
 buffer[303] = 8'h00;
 buffer[304] = 8'h00;
 buffer[305] = 8'h00;
 buffer[306] = 8'h66;
 buffer[307] = 8'h66;
 buffer[308] = 8'h66;
 buffer[309] = 8'h66;
 buffer[310] = 8'h66;
 buffer[311] = 8'h66;
 buffer[312] = 8'h66;
 buffer[313] = 8'h00;
 buffer[314] = 8'h66;
 buffer[315] = 8'h66;
 buffer[316] = 8'h00;
 buffer[317] = 8'h00;
 buffer[318] = 8'h00;
 buffer[319] = 8'h00;
 buffer[320] = 8'h00;
 buffer[321] = 8'h00;
 buffer[322] = 8'h7f;
 buffer[323] = 8'hdb;
 buffer[324] = 8'hdb;
 buffer[325] = 8'hdb;
 buffer[326] = 8'h7b;
 buffer[327] = 8'h1b;
 buffer[328] = 8'h1b;
 buffer[329] = 8'h1b;
 buffer[330] = 8'h1b;
 buffer[331] = 8'h1b;
 buffer[332] = 8'h00;
 buffer[333] = 8'h00;
 buffer[334] = 8'h00;
 buffer[335] = 8'h00;
 buffer[336] = 8'h00;
 buffer[337] = 8'h7c;
 buffer[338] = 8'hc6;
 buffer[339] = 8'h60;
 buffer[340] = 8'h38;
 buffer[341] = 8'h6c;
 buffer[342] = 8'hc6;
 buffer[343] = 8'hc6;
 buffer[344] = 8'h6c;
 buffer[345] = 8'h38;
 buffer[346] = 8'h0c;
 buffer[347] = 8'hc6;
 buffer[348] = 8'h7c;
 buffer[349] = 8'h00;
 buffer[350] = 8'h00;
 buffer[351] = 8'h00;
 buffer[352] = 8'h00;
 buffer[353] = 8'h00;
 buffer[354] = 8'h00;
 buffer[355] = 8'h00;
 buffer[356] = 8'h00;
 buffer[357] = 8'h00;
 buffer[358] = 8'h00;
 buffer[359] = 8'h00;
 buffer[360] = 8'hfe;
 buffer[361] = 8'hfe;
 buffer[362] = 8'hfe;
 buffer[363] = 8'hfe;
 buffer[364] = 8'h00;
 buffer[365] = 8'h00;
 buffer[366] = 8'h00;
 buffer[367] = 8'h00;
 buffer[368] = 8'h00;
 buffer[369] = 8'h00;
 buffer[370] = 8'h18;
 buffer[371] = 8'h3c;
 buffer[372] = 8'h7e;
 buffer[373] = 8'h18;
 buffer[374] = 8'h18;
 buffer[375] = 8'h18;
 buffer[376] = 8'h7e;
 buffer[377] = 8'h3c;
 buffer[378] = 8'h18;
 buffer[379] = 8'h7e;
 buffer[380] = 8'h00;
 buffer[381] = 8'h00;
 buffer[382] = 8'h00;
 buffer[383] = 8'h00;
 buffer[384] = 8'h00;
 buffer[385] = 8'h00;
 buffer[386] = 8'h18;
 buffer[387] = 8'h3c;
 buffer[388] = 8'h7e;
 buffer[389] = 8'h18;
 buffer[390] = 8'h18;
 buffer[391] = 8'h18;
 buffer[392] = 8'h18;
 buffer[393] = 8'h18;
 buffer[394] = 8'h18;
 buffer[395] = 8'h18;
 buffer[396] = 8'h00;
 buffer[397] = 8'h00;
 buffer[398] = 8'h00;
 buffer[399] = 8'h00;
 buffer[400] = 8'h00;
 buffer[401] = 8'h00;
 buffer[402] = 8'h18;
 buffer[403] = 8'h18;
 buffer[404] = 8'h18;
 buffer[405] = 8'h18;
 buffer[406] = 8'h18;
 buffer[407] = 8'h18;
 buffer[408] = 8'h18;
 buffer[409] = 8'h7e;
 buffer[410] = 8'h3c;
 buffer[411] = 8'h18;
 buffer[412] = 8'h00;
 buffer[413] = 8'h00;
 buffer[414] = 8'h00;
 buffer[415] = 8'h00;
 buffer[416] = 8'h00;
 buffer[417] = 8'h00;
 buffer[418] = 8'h00;
 buffer[419] = 8'h00;
 buffer[420] = 8'h00;
 buffer[421] = 8'h18;
 buffer[422] = 8'h0c;
 buffer[423] = 8'hfe;
 buffer[424] = 8'h0c;
 buffer[425] = 8'h18;
 buffer[426] = 8'h00;
 buffer[427] = 8'h00;
 buffer[428] = 8'h00;
 buffer[429] = 8'h00;
 buffer[430] = 8'h00;
 buffer[431] = 8'h00;
 buffer[432] = 8'h00;
 buffer[433] = 8'h00;
 buffer[434] = 8'h00;
 buffer[435] = 8'h00;
 buffer[436] = 8'h00;
 buffer[437] = 8'h30;
 buffer[438] = 8'h60;
 buffer[439] = 8'hfe;
 buffer[440] = 8'h60;
 buffer[441] = 8'h30;
 buffer[442] = 8'h00;
 buffer[443] = 8'h00;
 buffer[444] = 8'h00;
 buffer[445] = 8'h00;
 buffer[446] = 8'h00;
 buffer[447] = 8'h00;
 buffer[448] = 8'h00;
 buffer[449] = 8'h00;
 buffer[450] = 8'h00;
 buffer[451] = 8'h00;
 buffer[452] = 8'h00;
 buffer[453] = 8'h00;
 buffer[454] = 8'hc0;
 buffer[455] = 8'hc0;
 buffer[456] = 8'hc0;
 buffer[457] = 8'hfe;
 buffer[458] = 8'h00;
 buffer[459] = 8'h00;
 buffer[460] = 8'h00;
 buffer[461] = 8'h00;
 buffer[462] = 8'h00;
 buffer[463] = 8'h00;
 buffer[464] = 8'h00;
 buffer[465] = 8'h00;
 buffer[466] = 8'h00;
 buffer[467] = 8'h00;
 buffer[468] = 8'h00;
 buffer[469] = 8'h28;
 buffer[470] = 8'h6c;
 buffer[471] = 8'hfe;
 buffer[472] = 8'h6c;
 buffer[473] = 8'h28;
 buffer[474] = 8'h00;
 buffer[475] = 8'h00;
 buffer[476] = 8'h00;
 buffer[477] = 8'h00;
 buffer[478] = 8'h00;
 buffer[479] = 8'h00;
 buffer[480] = 8'h00;
 buffer[481] = 8'h00;
 buffer[482] = 8'h00;
 buffer[483] = 8'h00;
 buffer[484] = 8'h10;
 buffer[485] = 8'h38;
 buffer[486] = 8'h38;
 buffer[487] = 8'h7c;
 buffer[488] = 8'h7c;
 buffer[489] = 8'hfe;
 buffer[490] = 8'hfe;
 buffer[491] = 8'h00;
 buffer[492] = 8'h00;
 buffer[493] = 8'h00;
 buffer[494] = 8'h00;
 buffer[495] = 8'h00;
 buffer[496] = 8'h00;
 buffer[497] = 8'h00;
 buffer[498] = 8'h00;
 buffer[499] = 8'h00;
 buffer[500] = 8'hfe;
 buffer[501] = 8'hfe;
 buffer[502] = 8'h7c;
 buffer[503] = 8'h7c;
 buffer[504] = 8'h38;
 buffer[505] = 8'h38;
 buffer[506] = 8'h10;
 buffer[507] = 8'h00;
 buffer[508] = 8'h00;
 buffer[509] = 8'h00;
 buffer[510] = 8'h00;
 buffer[511] = 8'h00;
 buffer[512] = 8'h00;
 buffer[513] = 8'h00;
 buffer[514] = 8'h00;
 buffer[515] = 8'h00;
 buffer[516] = 8'h00;
 buffer[517] = 8'h00;
 buffer[518] = 8'h00;
 buffer[519] = 8'h00;
 buffer[520] = 8'h00;
 buffer[521] = 8'h00;
 buffer[522] = 8'h00;
 buffer[523] = 8'h00;
 buffer[524] = 8'h00;
 buffer[525] = 8'h00;
 buffer[526] = 8'h00;
 buffer[527] = 8'h00;
 buffer[528] = 8'h00;
 buffer[529] = 8'h00;
 buffer[530] = 8'h18;
 buffer[531] = 8'h3c;
 buffer[532] = 8'h3c;
 buffer[533] = 8'h3c;
 buffer[534] = 8'h18;
 buffer[535] = 8'h18;
 buffer[536] = 8'h18;
 buffer[537] = 8'h00;
 buffer[538] = 8'h18;
 buffer[539] = 8'h18;
 buffer[540] = 8'h00;
 buffer[541] = 8'h00;
 buffer[542] = 8'h00;
 buffer[543] = 8'h00;
 buffer[544] = 8'h00;
 buffer[545] = 8'h66;
 buffer[546] = 8'h66;
 buffer[547] = 8'h66;
 buffer[548] = 8'h24;
 buffer[549] = 8'h00;
 buffer[550] = 8'h00;
 buffer[551] = 8'h00;
 buffer[552] = 8'h00;
 buffer[553] = 8'h00;
 buffer[554] = 8'h00;
 buffer[555] = 8'h00;
 buffer[556] = 8'h00;
 buffer[557] = 8'h00;
 buffer[558] = 8'h00;
 buffer[559] = 8'h00;
 buffer[560] = 8'h00;
 buffer[561] = 8'h00;
 buffer[562] = 8'h00;
 buffer[563] = 8'h6c;
 buffer[564] = 8'h6c;
 buffer[565] = 8'hfe;
 buffer[566] = 8'h6c;
 buffer[567] = 8'h6c;
 buffer[568] = 8'h6c;
 buffer[569] = 8'hfe;
 buffer[570] = 8'h6c;
 buffer[571] = 8'h6c;
 buffer[572] = 8'h00;
 buffer[573] = 8'h00;
 buffer[574] = 8'h00;
 buffer[575] = 8'h00;
 buffer[576] = 8'h18;
 buffer[577] = 8'h18;
 buffer[578] = 8'h7c;
 buffer[579] = 8'hc6;
 buffer[580] = 8'hc2;
 buffer[581] = 8'hc0;
 buffer[582] = 8'h7c;
 buffer[583] = 8'h06;
 buffer[584] = 8'h06;
 buffer[585] = 8'h86;
 buffer[586] = 8'hc6;
 buffer[587] = 8'h7c;
 buffer[588] = 8'h18;
 buffer[589] = 8'h18;
 buffer[590] = 8'h00;
 buffer[591] = 8'h00;
 buffer[592] = 8'h00;
 buffer[593] = 8'h00;
 buffer[594] = 8'h00;
 buffer[595] = 8'h00;
 buffer[596] = 8'hc2;
 buffer[597] = 8'hc6;
 buffer[598] = 8'h0c;
 buffer[599] = 8'h18;
 buffer[600] = 8'h30;
 buffer[601] = 8'h60;
 buffer[602] = 8'hc6;
 buffer[603] = 8'h86;
 buffer[604] = 8'h00;
 buffer[605] = 8'h00;
 buffer[606] = 8'h00;
 buffer[607] = 8'h00;
 buffer[608] = 8'h00;
 buffer[609] = 8'h00;
 buffer[610] = 8'h38;
 buffer[611] = 8'h6c;
 buffer[612] = 8'h6c;
 buffer[613] = 8'h38;
 buffer[614] = 8'h76;
 buffer[615] = 8'hdc;
 buffer[616] = 8'hcc;
 buffer[617] = 8'hcc;
 buffer[618] = 8'hcc;
 buffer[619] = 8'h76;
 buffer[620] = 8'h00;
 buffer[621] = 8'h00;
 buffer[622] = 8'h00;
 buffer[623] = 8'h00;
 buffer[624] = 8'h00;
 buffer[625] = 8'h30;
 buffer[626] = 8'h30;
 buffer[627] = 8'h30;
 buffer[628] = 8'h60;
 buffer[629] = 8'h00;
 buffer[630] = 8'h00;
 buffer[631] = 8'h00;
 buffer[632] = 8'h00;
 buffer[633] = 8'h00;
 buffer[634] = 8'h00;
 buffer[635] = 8'h00;
 buffer[636] = 8'h00;
 buffer[637] = 8'h00;
 buffer[638] = 8'h00;
 buffer[639] = 8'h00;
 buffer[640] = 8'h00;
 buffer[641] = 8'h00;
 buffer[642] = 8'h0c;
 buffer[643] = 8'h18;
 buffer[644] = 8'h30;
 buffer[645] = 8'h30;
 buffer[646] = 8'h30;
 buffer[647] = 8'h30;
 buffer[648] = 8'h30;
 buffer[649] = 8'h30;
 buffer[650] = 8'h18;
 buffer[651] = 8'h0c;
 buffer[652] = 8'h00;
 buffer[653] = 8'h00;
 buffer[654] = 8'h00;
 buffer[655] = 8'h00;
 buffer[656] = 8'h00;
 buffer[657] = 8'h00;
 buffer[658] = 8'h30;
 buffer[659] = 8'h18;
 buffer[660] = 8'h0c;
 buffer[661] = 8'h0c;
 buffer[662] = 8'h0c;
 buffer[663] = 8'h0c;
 buffer[664] = 8'h0c;
 buffer[665] = 8'h0c;
 buffer[666] = 8'h18;
 buffer[667] = 8'h30;
 buffer[668] = 8'h00;
 buffer[669] = 8'h00;
 buffer[670] = 8'h00;
 buffer[671] = 8'h00;
 buffer[672] = 8'h00;
 buffer[673] = 8'h00;
 buffer[674] = 8'h00;
 buffer[675] = 8'h00;
 buffer[676] = 8'h00;
 buffer[677] = 8'h66;
 buffer[678] = 8'h3c;
 buffer[679] = 8'hff;
 buffer[680] = 8'h3c;
 buffer[681] = 8'h66;
 buffer[682] = 8'h00;
 buffer[683] = 8'h00;
 buffer[684] = 8'h00;
 buffer[685] = 8'h00;
 buffer[686] = 8'h00;
 buffer[687] = 8'h00;
 buffer[688] = 8'h00;
 buffer[689] = 8'h00;
 buffer[690] = 8'h00;
 buffer[691] = 8'h00;
 buffer[692] = 8'h00;
 buffer[693] = 8'h18;
 buffer[694] = 8'h18;
 buffer[695] = 8'h7e;
 buffer[696] = 8'h18;
 buffer[697] = 8'h18;
 buffer[698] = 8'h00;
 buffer[699] = 8'h00;
 buffer[700] = 8'h00;
 buffer[701] = 8'h00;
 buffer[702] = 8'h00;
 buffer[703] = 8'h00;
 buffer[704] = 8'h00;
 buffer[705] = 8'h00;
 buffer[706] = 8'h00;
 buffer[707] = 8'h00;
 buffer[708] = 8'h00;
 buffer[709] = 8'h00;
 buffer[710] = 8'h00;
 buffer[711] = 8'h00;
 buffer[712] = 8'h00;
 buffer[713] = 8'h18;
 buffer[714] = 8'h18;
 buffer[715] = 8'h18;
 buffer[716] = 8'h30;
 buffer[717] = 8'h00;
 buffer[718] = 8'h00;
 buffer[719] = 8'h00;
 buffer[720] = 8'h00;
 buffer[721] = 8'h00;
 buffer[722] = 8'h00;
 buffer[723] = 8'h00;
 buffer[724] = 8'h00;
 buffer[725] = 8'h00;
 buffer[726] = 8'h00;
 buffer[727] = 8'hfe;
 buffer[728] = 8'h00;
 buffer[729] = 8'h00;
 buffer[730] = 8'h00;
 buffer[731] = 8'h00;
 buffer[732] = 8'h00;
 buffer[733] = 8'h00;
 buffer[734] = 8'h00;
 buffer[735] = 8'h00;
 buffer[736] = 8'h00;
 buffer[737] = 8'h00;
 buffer[738] = 8'h00;
 buffer[739] = 8'h00;
 buffer[740] = 8'h00;
 buffer[741] = 8'h00;
 buffer[742] = 8'h00;
 buffer[743] = 8'h00;
 buffer[744] = 8'h00;
 buffer[745] = 8'h00;
 buffer[746] = 8'h18;
 buffer[747] = 8'h18;
 buffer[748] = 8'h00;
 buffer[749] = 8'h00;
 buffer[750] = 8'h00;
 buffer[751] = 8'h00;
 buffer[752] = 8'h00;
 buffer[753] = 8'h00;
 buffer[754] = 8'h00;
 buffer[755] = 8'h00;
 buffer[756] = 8'h02;
 buffer[757] = 8'h06;
 buffer[758] = 8'h0c;
 buffer[759] = 8'h18;
 buffer[760] = 8'h30;
 buffer[761] = 8'h60;
 buffer[762] = 8'hc0;
 buffer[763] = 8'h80;
 buffer[764] = 8'h00;
 buffer[765] = 8'h00;
 buffer[766] = 8'h00;
 buffer[767] = 8'h00;
 buffer[768] = 8'h00;
 buffer[769] = 8'h00;
 buffer[770] = 8'h38;
 buffer[771] = 8'h6c;
 buffer[772] = 8'hc6;
 buffer[773] = 8'hc6;
 buffer[774] = 8'hd6;
 buffer[775] = 8'hd6;
 buffer[776] = 8'hc6;
 buffer[777] = 8'hc6;
 buffer[778] = 8'h6c;
 buffer[779] = 8'h38;
 buffer[780] = 8'h00;
 buffer[781] = 8'h00;
 buffer[782] = 8'h00;
 buffer[783] = 8'h00;
 buffer[784] = 8'h00;
 buffer[785] = 8'h00;
 buffer[786] = 8'h18;
 buffer[787] = 8'h38;
 buffer[788] = 8'h78;
 buffer[789] = 8'h18;
 buffer[790] = 8'h18;
 buffer[791] = 8'h18;
 buffer[792] = 8'h18;
 buffer[793] = 8'h18;
 buffer[794] = 8'h18;
 buffer[795] = 8'h7e;
 buffer[796] = 8'h00;
 buffer[797] = 8'h00;
 buffer[798] = 8'h00;
 buffer[799] = 8'h00;
 buffer[800] = 8'h00;
 buffer[801] = 8'h00;
 buffer[802] = 8'h7c;
 buffer[803] = 8'hc6;
 buffer[804] = 8'h06;
 buffer[805] = 8'h0c;
 buffer[806] = 8'h18;
 buffer[807] = 8'h30;
 buffer[808] = 8'h60;
 buffer[809] = 8'hc0;
 buffer[810] = 8'hc6;
 buffer[811] = 8'hfe;
 buffer[812] = 8'h00;
 buffer[813] = 8'h00;
 buffer[814] = 8'h00;
 buffer[815] = 8'h00;
 buffer[816] = 8'h00;
 buffer[817] = 8'h00;
 buffer[818] = 8'h7c;
 buffer[819] = 8'hc6;
 buffer[820] = 8'h06;
 buffer[821] = 8'h06;
 buffer[822] = 8'h3c;
 buffer[823] = 8'h06;
 buffer[824] = 8'h06;
 buffer[825] = 8'h06;
 buffer[826] = 8'hc6;
 buffer[827] = 8'h7c;
 buffer[828] = 8'h00;
 buffer[829] = 8'h00;
 buffer[830] = 8'h00;
 buffer[831] = 8'h00;
 buffer[832] = 8'h00;
 buffer[833] = 8'h00;
 buffer[834] = 8'h0c;
 buffer[835] = 8'h1c;
 buffer[836] = 8'h3c;
 buffer[837] = 8'h6c;
 buffer[838] = 8'hcc;
 buffer[839] = 8'hfe;
 buffer[840] = 8'h0c;
 buffer[841] = 8'h0c;
 buffer[842] = 8'h0c;
 buffer[843] = 8'h1e;
 buffer[844] = 8'h00;
 buffer[845] = 8'h00;
 buffer[846] = 8'h00;
 buffer[847] = 8'h00;
 buffer[848] = 8'h00;
 buffer[849] = 8'h00;
 buffer[850] = 8'hfe;
 buffer[851] = 8'hc0;
 buffer[852] = 8'hc0;
 buffer[853] = 8'hc0;
 buffer[854] = 8'hfc;
 buffer[855] = 8'h06;
 buffer[856] = 8'h06;
 buffer[857] = 8'h06;
 buffer[858] = 8'hc6;
 buffer[859] = 8'h7c;
 buffer[860] = 8'h00;
 buffer[861] = 8'h00;
 buffer[862] = 8'h00;
 buffer[863] = 8'h00;
 buffer[864] = 8'h00;
 buffer[865] = 8'h00;
 buffer[866] = 8'h38;
 buffer[867] = 8'h60;
 buffer[868] = 8'hc0;
 buffer[869] = 8'hc0;
 buffer[870] = 8'hfc;
 buffer[871] = 8'hc6;
 buffer[872] = 8'hc6;
 buffer[873] = 8'hc6;
 buffer[874] = 8'hc6;
 buffer[875] = 8'h7c;
 buffer[876] = 8'h00;
 buffer[877] = 8'h00;
 buffer[878] = 8'h00;
 buffer[879] = 8'h00;
 buffer[880] = 8'h00;
 buffer[881] = 8'h00;
 buffer[882] = 8'hfe;
 buffer[883] = 8'hc6;
 buffer[884] = 8'h06;
 buffer[885] = 8'h06;
 buffer[886] = 8'h0c;
 buffer[887] = 8'h18;
 buffer[888] = 8'h30;
 buffer[889] = 8'h30;
 buffer[890] = 8'h30;
 buffer[891] = 8'h30;
 buffer[892] = 8'h00;
 buffer[893] = 8'h00;
 buffer[894] = 8'h00;
 buffer[895] = 8'h00;
 buffer[896] = 8'h00;
 buffer[897] = 8'h00;
 buffer[898] = 8'h7c;
 buffer[899] = 8'hc6;
 buffer[900] = 8'hc6;
 buffer[901] = 8'hc6;
 buffer[902] = 8'h7c;
 buffer[903] = 8'hc6;
 buffer[904] = 8'hc6;
 buffer[905] = 8'hc6;
 buffer[906] = 8'hc6;
 buffer[907] = 8'h7c;
 buffer[908] = 8'h00;
 buffer[909] = 8'h00;
 buffer[910] = 8'h00;
 buffer[911] = 8'h00;
 buffer[912] = 8'h00;
 buffer[913] = 8'h00;
 buffer[914] = 8'h7c;
 buffer[915] = 8'hc6;
 buffer[916] = 8'hc6;
 buffer[917] = 8'hc6;
 buffer[918] = 8'h7e;
 buffer[919] = 8'h06;
 buffer[920] = 8'h06;
 buffer[921] = 8'h06;
 buffer[922] = 8'h0c;
 buffer[923] = 8'h78;
 buffer[924] = 8'h00;
 buffer[925] = 8'h00;
 buffer[926] = 8'h00;
 buffer[927] = 8'h00;
 buffer[928] = 8'h00;
 buffer[929] = 8'h00;
 buffer[930] = 8'h00;
 buffer[931] = 8'h00;
 buffer[932] = 8'h18;
 buffer[933] = 8'h18;
 buffer[934] = 8'h00;
 buffer[935] = 8'h00;
 buffer[936] = 8'h00;
 buffer[937] = 8'h18;
 buffer[938] = 8'h18;
 buffer[939] = 8'h00;
 buffer[940] = 8'h00;
 buffer[941] = 8'h00;
 buffer[942] = 8'h00;
 buffer[943] = 8'h00;
 buffer[944] = 8'h00;
 buffer[945] = 8'h00;
 buffer[946] = 8'h00;
 buffer[947] = 8'h00;
 buffer[948] = 8'h18;
 buffer[949] = 8'h18;
 buffer[950] = 8'h00;
 buffer[951] = 8'h00;
 buffer[952] = 8'h00;
 buffer[953] = 8'h18;
 buffer[954] = 8'h18;
 buffer[955] = 8'h30;
 buffer[956] = 8'h00;
 buffer[957] = 8'h00;
 buffer[958] = 8'h00;
 buffer[959] = 8'h00;
 buffer[960] = 8'h00;
 buffer[961] = 8'h00;
 buffer[962] = 8'h00;
 buffer[963] = 8'h06;
 buffer[964] = 8'h0c;
 buffer[965] = 8'h18;
 buffer[966] = 8'h30;
 buffer[967] = 8'h60;
 buffer[968] = 8'h30;
 buffer[969] = 8'h18;
 buffer[970] = 8'h0c;
 buffer[971] = 8'h06;
 buffer[972] = 8'h00;
 buffer[973] = 8'h00;
 buffer[974] = 8'h00;
 buffer[975] = 8'h00;
 buffer[976] = 8'h00;
 buffer[977] = 8'h00;
 buffer[978] = 8'h00;
 buffer[979] = 8'h00;
 buffer[980] = 8'h00;
 buffer[981] = 8'h7e;
 buffer[982] = 8'h00;
 buffer[983] = 8'h00;
 buffer[984] = 8'h7e;
 buffer[985] = 8'h00;
 buffer[986] = 8'h00;
 buffer[987] = 8'h00;
 buffer[988] = 8'h00;
 buffer[989] = 8'h00;
 buffer[990] = 8'h00;
 buffer[991] = 8'h00;
 buffer[992] = 8'h00;
 buffer[993] = 8'h00;
 buffer[994] = 8'h00;
 buffer[995] = 8'h60;
 buffer[996] = 8'h30;
 buffer[997] = 8'h18;
 buffer[998] = 8'h0c;
 buffer[999] = 8'h06;
 buffer[1000] = 8'h0c;
 buffer[1001] = 8'h18;
 buffer[1002] = 8'h30;
 buffer[1003] = 8'h60;
 buffer[1004] = 8'h00;
 buffer[1005] = 8'h00;
 buffer[1006] = 8'h00;
 buffer[1007] = 8'h00;
 buffer[1008] = 8'h00;
 buffer[1009] = 8'h00;
 buffer[1010] = 8'h7c;
 buffer[1011] = 8'hc6;
 buffer[1012] = 8'hc6;
 buffer[1013] = 8'h0c;
 buffer[1014] = 8'h18;
 buffer[1015] = 8'h18;
 buffer[1016] = 8'h18;
 buffer[1017] = 8'h00;
 buffer[1018] = 8'h18;
 buffer[1019] = 8'h18;
 buffer[1020] = 8'h00;
 buffer[1021] = 8'h00;
 buffer[1022] = 8'h00;
 buffer[1023] = 8'h00;
 buffer[1024] = 8'h00;
 buffer[1025] = 8'h00;
 buffer[1026] = 8'h00;
 buffer[1027] = 8'h7c;
 buffer[1028] = 8'hc6;
 buffer[1029] = 8'hc6;
 buffer[1030] = 8'hde;
 buffer[1031] = 8'hde;
 buffer[1032] = 8'hde;
 buffer[1033] = 8'hdc;
 buffer[1034] = 8'hc0;
 buffer[1035] = 8'h7c;
 buffer[1036] = 8'h00;
 buffer[1037] = 8'h00;
 buffer[1038] = 8'h00;
 buffer[1039] = 8'h00;
 buffer[1040] = 8'h00;
 buffer[1041] = 8'h00;
 buffer[1042] = 8'h10;
 buffer[1043] = 8'h38;
 buffer[1044] = 8'h6c;
 buffer[1045] = 8'hc6;
 buffer[1046] = 8'hc6;
 buffer[1047] = 8'hfe;
 buffer[1048] = 8'hc6;
 buffer[1049] = 8'hc6;
 buffer[1050] = 8'hc6;
 buffer[1051] = 8'hc6;
 buffer[1052] = 8'h00;
 buffer[1053] = 8'h00;
 buffer[1054] = 8'h00;
 buffer[1055] = 8'h00;
 buffer[1056] = 8'h00;
 buffer[1057] = 8'h00;
 buffer[1058] = 8'hfc;
 buffer[1059] = 8'h66;
 buffer[1060] = 8'h66;
 buffer[1061] = 8'h66;
 buffer[1062] = 8'h7c;
 buffer[1063] = 8'h66;
 buffer[1064] = 8'h66;
 buffer[1065] = 8'h66;
 buffer[1066] = 8'h66;
 buffer[1067] = 8'hfc;
 buffer[1068] = 8'h00;
 buffer[1069] = 8'h00;
 buffer[1070] = 8'h00;
 buffer[1071] = 8'h00;
 buffer[1072] = 8'h00;
 buffer[1073] = 8'h00;
 buffer[1074] = 8'h3c;
 buffer[1075] = 8'h66;
 buffer[1076] = 8'hc2;
 buffer[1077] = 8'hc0;
 buffer[1078] = 8'hc0;
 buffer[1079] = 8'hc0;
 buffer[1080] = 8'hc0;
 buffer[1081] = 8'hc2;
 buffer[1082] = 8'h66;
 buffer[1083] = 8'h3c;
 buffer[1084] = 8'h00;
 buffer[1085] = 8'h00;
 buffer[1086] = 8'h00;
 buffer[1087] = 8'h00;
 buffer[1088] = 8'h00;
 buffer[1089] = 8'h00;
 buffer[1090] = 8'hf8;
 buffer[1091] = 8'h6c;
 buffer[1092] = 8'h66;
 buffer[1093] = 8'h66;
 buffer[1094] = 8'h66;
 buffer[1095] = 8'h66;
 buffer[1096] = 8'h66;
 buffer[1097] = 8'h66;
 buffer[1098] = 8'h6c;
 buffer[1099] = 8'hf8;
 buffer[1100] = 8'h00;
 buffer[1101] = 8'h00;
 buffer[1102] = 8'h00;
 buffer[1103] = 8'h00;
 buffer[1104] = 8'h00;
 buffer[1105] = 8'h00;
 buffer[1106] = 8'hfe;
 buffer[1107] = 8'h66;
 buffer[1108] = 8'h62;
 buffer[1109] = 8'h68;
 buffer[1110] = 8'h78;
 buffer[1111] = 8'h68;
 buffer[1112] = 8'h60;
 buffer[1113] = 8'h62;
 buffer[1114] = 8'h66;
 buffer[1115] = 8'hfe;
 buffer[1116] = 8'h00;
 buffer[1117] = 8'h00;
 buffer[1118] = 8'h00;
 buffer[1119] = 8'h00;
 buffer[1120] = 8'h00;
 buffer[1121] = 8'h00;
 buffer[1122] = 8'hfe;
 buffer[1123] = 8'h66;
 buffer[1124] = 8'h62;
 buffer[1125] = 8'h68;
 buffer[1126] = 8'h78;
 buffer[1127] = 8'h68;
 buffer[1128] = 8'h60;
 buffer[1129] = 8'h60;
 buffer[1130] = 8'h60;
 buffer[1131] = 8'hf0;
 buffer[1132] = 8'h00;
 buffer[1133] = 8'h00;
 buffer[1134] = 8'h00;
 buffer[1135] = 8'h00;
 buffer[1136] = 8'h00;
 buffer[1137] = 8'h00;
 buffer[1138] = 8'h3c;
 buffer[1139] = 8'h66;
 buffer[1140] = 8'hc2;
 buffer[1141] = 8'hc0;
 buffer[1142] = 8'hc0;
 buffer[1143] = 8'hde;
 buffer[1144] = 8'hc6;
 buffer[1145] = 8'hc6;
 buffer[1146] = 8'h66;
 buffer[1147] = 8'h3a;
 buffer[1148] = 8'h00;
 buffer[1149] = 8'h00;
 buffer[1150] = 8'h00;
 buffer[1151] = 8'h00;
 buffer[1152] = 8'h00;
 buffer[1153] = 8'h00;
 buffer[1154] = 8'hc6;
 buffer[1155] = 8'hc6;
 buffer[1156] = 8'hc6;
 buffer[1157] = 8'hc6;
 buffer[1158] = 8'hfe;
 buffer[1159] = 8'hc6;
 buffer[1160] = 8'hc6;
 buffer[1161] = 8'hc6;
 buffer[1162] = 8'hc6;
 buffer[1163] = 8'hc6;
 buffer[1164] = 8'h00;
 buffer[1165] = 8'h00;
 buffer[1166] = 8'h00;
 buffer[1167] = 8'h00;
 buffer[1168] = 8'h00;
 buffer[1169] = 8'h00;
 buffer[1170] = 8'h3c;
 buffer[1171] = 8'h18;
 buffer[1172] = 8'h18;
 buffer[1173] = 8'h18;
 buffer[1174] = 8'h18;
 buffer[1175] = 8'h18;
 buffer[1176] = 8'h18;
 buffer[1177] = 8'h18;
 buffer[1178] = 8'h18;
 buffer[1179] = 8'h3c;
 buffer[1180] = 8'h00;
 buffer[1181] = 8'h00;
 buffer[1182] = 8'h00;
 buffer[1183] = 8'h00;
 buffer[1184] = 8'h00;
 buffer[1185] = 8'h00;
 buffer[1186] = 8'h1e;
 buffer[1187] = 8'h0c;
 buffer[1188] = 8'h0c;
 buffer[1189] = 8'h0c;
 buffer[1190] = 8'h0c;
 buffer[1191] = 8'h0c;
 buffer[1192] = 8'hcc;
 buffer[1193] = 8'hcc;
 buffer[1194] = 8'hcc;
 buffer[1195] = 8'h78;
 buffer[1196] = 8'h00;
 buffer[1197] = 8'h00;
 buffer[1198] = 8'h00;
 buffer[1199] = 8'h00;
 buffer[1200] = 8'h00;
 buffer[1201] = 8'h00;
 buffer[1202] = 8'he6;
 buffer[1203] = 8'h66;
 buffer[1204] = 8'h66;
 buffer[1205] = 8'h6c;
 buffer[1206] = 8'h78;
 buffer[1207] = 8'h78;
 buffer[1208] = 8'h6c;
 buffer[1209] = 8'h66;
 buffer[1210] = 8'h66;
 buffer[1211] = 8'he6;
 buffer[1212] = 8'h00;
 buffer[1213] = 8'h00;
 buffer[1214] = 8'h00;
 buffer[1215] = 8'h00;
 buffer[1216] = 8'h00;
 buffer[1217] = 8'h00;
 buffer[1218] = 8'hf0;
 buffer[1219] = 8'h60;
 buffer[1220] = 8'h60;
 buffer[1221] = 8'h60;
 buffer[1222] = 8'h60;
 buffer[1223] = 8'h60;
 buffer[1224] = 8'h60;
 buffer[1225] = 8'h62;
 buffer[1226] = 8'h66;
 buffer[1227] = 8'hfe;
 buffer[1228] = 8'h00;
 buffer[1229] = 8'h00;
 buffer[1230] = 8'h00;
 buffer[1231] = 8'h00;
 buffer[1232] = 8'h00;
 buffer[1233] = 8'h00;
 buffer[1234] = 8'hc6;
 buffer[1235] = 8'hee;
 buffer[1236] = 8'hfe;
 buffer[1237] = 8'hfe;
 buffer[1238] = 8'hd6;
 buffer[1239] = 8'hc6;
 buffer[1240] = 8'hc6;
 buffer[1241] = 8'hc6;
 buffer[1242] = 8'hc6;
 buffer[1243] = 8'hc6;
 buffer[1244] = 8'h00;
 buffer[1245] = 8'h00;
 buffer[1246] = 8'h00;
 buffer[1247] = 8'h00;
 buffer[1248] = 8'h00;
 buffer[1249] = 8'h00;
 buffer[1250] = 8'hc6;
 buffer[1251] = 8'he6;
 buffer[1252] = 8'hf6;
 buffer[1253] = 8'hfe;
 buffer[1254] = 8'hde;
 buffer[1255] = 8'hce;
 buffer[1256] = 8'hc6;
 buffer[1257] = 8'hc6;
 buffer[1258] = 8'hc6;
 buffer[1259] = 8'hc6;
 buffer[1260] = 8'h00;
 buffer[1261] = 8'h00;
 buffer[1262] = 8'h00;
 buffer[1263] = 8'h00;
 buffer[1264] = 8'h00;
 buffer[1265] = 8'h00;
 buffer[1266] = 8'h7c;
 buffer[1267] = 8'hc6;
 buffer[1268] = 8'hc6;
 buffer[1269] = 8'hc6;
 buffer[1270] = 8'hc6;
 buffer[1271] = 8'hc6;
 buffer[1272] = 8'hc6;
 buffer[1273] = 8'hc6;
 buffer[1274] = 8'hc6;
 buffer[1275] = 8'h7c;
 buffer[1276] = 8'h00;
 buffer[1277] = 8'h00;
 buffer[1278] = 8'h00;
 buffer[1279] = 8'h00;
 buffer[1280] = 8'h00;
 buffer[1281] = 8'h00;
 buffer[1282] = 8'hfc;
 buffer[1283] = 8'h66;
 buffer[1284] = 8'h66;
 buffer[1285] = 8'h66;
 buffer[1286] = 8'h7c;
 buffer[1287] = 8'h60;
 buffer[1288] = 8'h60;
 buffer[1289] = 8'h60;
 buffer[1290] = 8'h60;
 buffer[1291] = 8'hf0;
 buffer[1292] = 8'h00;
 buffer[1293] = 8'h00;
 buffer[1294] = 8'h00;
 buffer[1295] = 8'h00;
 buffer[1296] = 8'h00;
 buffer[1297] = 8'h00;
 buffer[1298] = 8'h7c;
 buffer[1299] = 8'hc6;
 buffer[1300] = 8'hc6;
 buffer[1301] = 8'hc6;
 buffer[1302] = 8'hc6;
 buffer[1303] = 8'hc6;
 buffer[1304] = 8'hc6;
 buffer[1305] = 8'hd6;
 buffer[1306] = 8'hde;
 buffer[1307] = 8'h7c;
 buffer[1308] = 8'h0c;
 buffer[1309] = 8'h0e;
 buffer[1310] = 8'h00;
 buffer[1311] = 8'h00;
 buffer[1312] = 8'h00;
 buffer[1313] = 8'h00;
 buffer[1314] = 8'hfc;
 buffer[1315] = 8'h66;
 buffer[1316] = 8'h66;
 buffer[1317] = 8'h66;
 buffer[1318] = 8'h7c;
 buffer[1319] = 8'h6c;
 buffer[1320] = 8'h66;
 buffer[1321] = 8'h66;
 buffer[1322] = 8'h66;
 buffer[1323] = 8'he6;
 buffer[1324] = 8'h00;
 buffer[1325] = 8'h00;
 buffer[1326] = 8'h00;
 buffer[1327] = 8'h00;
 buffer[1328] = 8'h00;
 buffer[1329] = 8'h00;
 buffer[1330] = 8'h7c;
 buffer[1331] = 8'hc6;
 buffer[1332] = 8'hc6;
 buffer[1333] = 8'h60;
 buffer[1334] = 8'h38;
 buffer[1335] = 8'h0c;
 buffer[1336] = 8'h06;
 buffer[1337] = 8'hc6;
 buffer[1338] = 8'hc6;
 buffer[1339] = 8'h7c;
 buffer[1340] = 8'h00;
 buffer[1341] = 8'h00;
 buffer[1342] = 8'h00;
 buffer[1343] = 8'h00;
 buffer[1344] = 8'h00;
 buffer[1345] = 8'h00;
 buffer[1346] = 8'h7e;
 buffer[1347] = 8'h7e;
 buffer[1348] = 8'h5a;
 buffer[1349] = 8'h18;
 buffer[1350] = 8'h18;
 buffer[1351] = 8'h18;
 buffer[1352] = 8'h18;
 buffer[1353] = 8'h18;
 buffer[1354] = 8'h18;
 buffer[1355] = 8'h3c;
 buffer[1356] = 8'h00;
 buffer[1357] = 8'h00;
 buffer[1358] = 8'h00;
 buffer[1359] = 8'h00;
 buffer[1360] = 8'h00;
 buffer[1361] = 8'h00;
 buffer[1362] = 8'hc6;
 buffer[1363] = 8'hc6;
 buffer[1364] = 8'hc6;
 buffer[1365] = 8'hc6;
 buffer[1366] = 8'hc6;
 buffer[1367] = 8'hc6;
 buffer[1368] = 8'hc6;
 buffer[1369] = 8'hc6;
 buffer[1370] = 8'hc6;
 buffer[1371] = 8'h7c;
 buffer[1372] = 8'h00;
 buffer[1373] = 8'h00;
 buffer[1374] = 8'h00;
 buffer[1375] = 8'h00;
 buffer[1376] = 8'h00;
 buffer[1377] = 8'h00;
 buffer[1378] = 8'hc6;
 buffer[1379] = 8'hc6;
 buffer[1380] = 8'hc6;
 buffer[1381] = 8'hc6;
 buffer[1382] = 8'hc6;
 buffer[1383] = 8'hc6;
 buffer[1384] = 8'hc6;
 buffer[1385] = 8'h6c;
 buffer[1386] = 8'h38;
 buffer[1387] = 8'h10;
 buffer[1388] = 8'h00;
 buffer[1389] = 8'h00;
 buffer[1390] = 8'h00;
 buffer[1391] = 8'h00;
 buffer[1392] = 8'h00;
 buffer[1393] = 8'h00;
 buffer[1394] = 8'hc6;
 buffer[1395] = 8'hc6;
 buffer[1396] = 8'hc6;
 buffer[1397] = 8'hc6;
 buffer[1398] = 8'hd6;
 buffer[1399] = 8'hd6;
 buffer[1400] = 8'hd6;
 buffer[1401] = 8'hfe;
 buffer[1402] = 8'hee;
 buffer[1403] = 8'h6c;
 buffer[1404] = 8'h00;
 buffer[1405] = 8'h00;
 buffer[1406] = 8'h00;
 buffer[1407] = 8'h00;
 buffer[1408] = 8'h00;
 buffer[1409] = 8'h00;
 buffer[1410] = 8'hc6;
 buffer[1411] = 8'hc6;
 buffer[1412] = 8'h6c;
 buffer[1413] = 8'h7c;
 buffer[1414] = 8'h38;
 buffer[1415] = 8'h38;
 buffer[1416] = 8'h7c;
 buffer[1417] = 8'h6c;
 buffer[1418] = 8'hc6;
 buffer[1419] = 8'hc6;
 buffer[1420] = 8'h00;
 buffer[1421] = 8'h00;
 buffer[1422] = 8'h00;
 buffer[1423] = 8'h00;
 buffer[1424] = 8'h00;
 buffer[1425] = 8'h00;
 buffer[1426] = 8'h66;
 buffer[1427] = 8'h66;
 buffer[1428] = 8'h66;
 buffer[1429] = 8'h66;
 buffer[1430] = 8'h3c;
 buffer[1431] = 8'h18;
 buffer[1432] = 8'h18;
 buffer[1433] = 8'h18;
 buffer[1434] = 8'h18;
 buffer[1435] = 8'h3c;
 buffer[1436] = 8'h00;
 buffer[1437] = 8'h00;
 buffer[1438] = 8'h00;
 buffer[1439] = 8'h00;
 buffer[1440] = 8'h00;
 buffer[1441] = 8'h00;
 buffer[1442] = 8'hfe;
 buffer[1443] = 8'hc6;
 buffer[1444] = 8'h86;
 buffer[1445] = 8'h0c;
 buffer[1446] = 8'h18;
 buffer[1447] = 8'h30;
 buffer[1448] = 8'h60;
 buffer[1449] = 8'hc2;
 buffer[1450] = 8'hc6;
 buffer[1451] = 8'hfe;
 buffer[1452] = 8'h00;
 buffer[1453] = 8'h00;
 buffer[1454] = 8'h00;
 buffer[1455] = 8'h00;
 buffer[1456] = 8'h00;
 buffer[1457] = 8'h00;
 buffer[1458] = 8'h3c;
 buffer[1459] = 8'h30;
 buffer[1460] = 8'h30;
 buffer[1461] = 8'h30;
 buffer[1462] = 8'h30;
 buffer[1463] = 8'h30;
 buffer[1464] = 8'h30;
 buffer[1465] = 8'h30;
 buffer[1466] = 8'h30;
 buffer[1467] = 8'h3c;
 buffer[1468] = 8'h00;
 buffer[1469] = 8'h00;
 buffer[1470] = 8'h00;
 buffer[1471] = 8'h00;
 buffer[1472] = 8'h00;
 buffer[1473] = 8'h00;
 buffer[1474] = 8'h00;
 buffer[1475] = 8'h80;
 buffer[1476] = 8'hc0;
 buffer[1477] = 8'he0;
 buffer[1478] = 8'h70;
 buffer[1479] = 8'h38;
 buffer[1480] = 8'h1c;
 buffer[1481] = 8'h0e;
 buffer[1482] = 8'h06;
 buffer[1483] = 8'h02;
 buffer[1484] = 8'h00;
 buffer[1485] = 8'h00;
 buffer[1486] = 8'h00;
 buffer[1487] = 8'h00;
 buffer[1488] = 8'h00;
 buffer[1489] = 8'h00;
 buffer[1490] = 8'h3c;
 buffer[1491] = 8'h0c;
 buffer[1492] = 8'h0c;
 buffer[1493] = 8'h0c;
 buffer[1494] = 8'h0c;
 buffer[1495] = 8'h0c;
 buffer[1496] = 8'h0c;
 buffer[1497] = 8'h0c;
 buffer[1498] = 8'h0c;
 buffer[1499] = 8'h3c;
 buffer[1500] = 8'h00;
 buffer[1501] = 8'h00;
 buffer[1502] = 8'h00;
 buffer[1503] = 8'h00;
 buffer[1504] = 8'h10;
 buffer[1505] = 8'h38;
 buffer[1506] = 8'h6c;
 buffer[1507] = 8'hc6;
 buffer[1508] = 8'h00;
 buffer[1509] = 8'h00;
 buffer[1510] = 8'h00;
 buffer[1511] = 8'h00;
 buffer[1512] = 8'h00;
 buffer[1513] = 8'h00;
 buffer[1514] = 8'h00;
 buffer[1515] = 8'h00;
 buffer[1516] = 8'h00;
 buffer[1517] = 8'h00;
 buffer[1518] = 8'h00;
 buffer[1519] = 8'h00;
 buffer[1520] = 8'h00;
 buffer[1521] = 8'h00;
 buffer[1522] = 8'h00;
 buffer[1523] = 8'h00;
 buffer[1524] = 8'h00;
 buffer[1525] = 8'h00;
 buffer[1526] = 8'h00;
 buffer[1527] = 8'h00;
 buffer[1528] = 8'h00;
 buffer[1529] = 8'h00;
 buffer[1530] = 8'h00;
 buffer[1531] = 8'h00;
 buffer[1532] = 8'h00;
 buffer[1533] = 8'hff;
 buffer[1534] = 8'h00;
 buffer[1535] = 8'h00;
 buffer[1536] = 8'h30;
 buffer[1537] = 8'h30;
 buffer[1538] = 8'h18;
 buffer[1539] = 8'h00;
 buffer[1540] = 8'h00;
 buffer[1541] = 8'h00;
 buffer[1542] = 8'h00;
 buffer[1543] = 8'h00;
 buffer[1544] = 8'h00;
 buffer[1545] = 8'h00;
 buffer[1546] = 8'h00;
 buffer[1547] = 8'h00;
 buffer[1548] = 8'h00;
 buffer[1549] = 8'h00;
 buffer[1550] = 8'h00;
 buffer[1551] = 8'h00;
 buffer[1552] = 8'h00;
 buffer[1553] = 8'h00;
 buffer[1554] = 8'h00;
 buffer[1555] = 8'h00;
 buffer[1556] = 8'h00;
 buffer[1557] = 8'h78;
 buffer[1558] = 8'h0c;
 buffer[1559] = 8'h7c;
 buffer[1560] = 8'hcc;
 buffer[1561] = 8'hcc;
 buffer[1562] = 8'hcc;
 buffer[1563] = 8'h76;
 buffer[1564] = 8'h00;
 buffer[1565] = 8'h00;
 buffer[1566] = 8'h00;
 buffer[1567] = 8'h00;
 buffer[1568] = 8'h00;
 buffer[1569] = 8'h00;
 buffer[1570] = 8'he0;
 buffer[1571] = 8'h60;
 buffer[1572] = 8'h60;
 buffer[1573] = 8'h78;
 buffer[1574] = 8'h6c;
 buffer[1575] = 8'h66;
 buffer[1576] = 8'h66;
 buffer[1577] = 8'h66;
 buffer[1578] = 8'h66;
 buffer[1579] = 8'h7c;
 buffer[1580] = 8'h00;
 buffer[1581] = 8'h00;
 buffer[1582] = 8'h00;
 buffer[1583] = 8'h00;
 buffer[1584] = 8'h00;
 buffer[1585] = 8'h00;
 buffer[1586] = 8'h00;
 buffer[1587] = 8'h00;
 buffer[1588] = 8'h00;
 buffer[1589] = 8'h7c;
 buffer[1590] = 8'hc6;
 buffer[1591] = 8'hc0;
 buffer[1592] = 8'hc0;
 buffer[1593] = 8'hc0;
 buffer[1594] = 8'hc6;
 buffer[1595] = 8'h7c;
 buffer[1596] = 8'h00;
 buffer[1597] = 8'h00;
 buffer[1598] = 8'h00;
 buffer[1599] = 8'h00;
 buffer[1600] = 8'h00;
 buffer[1601] = 8'h00;
 buffer[1602] = 8'h1c;
 buffer[1603] = 8'h0c;
 buffer[1604] = 8'h0c;
 buffer[1605] = 8'h3c;
 buffer[1606] = 8'h6c;
 buffer[1607] = 8'hcc;
 buffer[1608] = 8'hcc;
 buffer[1609] = 8'hcc;
 buffer[1610] = 8'hcc;
 buffer[1611] = 8'h76;
 buffer[1612] = 8'h00;
 buffer[1613] = 8'h00;
 buffer[1614] = 8'h00;
 buffer[1615] = 8'h00;
 buffer[1616] = 8'h00;
 buffer[1617] = 8'h00;
 buffer[1618] = 8'h00;
 buffer[1619] = 8'h00;
 buffer[1620] = 8'h00;
 buffer[1621] = 8'h7c;
 buffer[1622] = 8'hc6;
 buffer[1623] = 8'hfe;
 buffer[1624] = 8'hc0;
 buffer[1625] = 8'hc0;
 buffer[1626] = 8'hc6;
 buffer[1627] = 8'h7c;
 buffer[1628] = 8'h00;
 buffer[1629] = 8'h00;
 buffer[1630] = 8'h00;
 buffer[1631] = 8'h00;
 buffer[1632] = 8'h00;
 buffer[1633] = 8'h00;
 buffer[1634] = 8'h38;
 buffer[1635] = 8'h6c;
 buffer[1636] = 8'h64;
 buffer[1637] = 8'h60;
 buffer[1638] = 8'hf0;
 buffer[1639] = 8'h60;
 buffer[1640] = 8'h60;
 buffer[1641] = 8'h60;
 buffer[1642] = 8'h60;
 buffer[1643] = 8'hf0;
 buffer[1644] = 8'h00;
 buffer[1645] = 8'h00;
 buffer[1646] = 8'h00;
 buffer[1647] = 8'h00;
 buffer[1648] = 8'h00;
 buffer[1649] = 8'h00;
 buffer[1650] = 8'h00;
 buffer[1651] = 8'h00;
 buffer[1652] = 8'h00;
 buffer[1653] = 8'h76;
 buffer[1654] = 8'hcc;
 buffer[1655] = 8'hcc;
 buffer[1656] = 8'hcc;
 buffer[1657] = 8'hcc;
 buffer[1658] = 8'hcc;
 buffer[1659] = 8'h7c;
 buffer[1660] = 8'h0c;
 buffer[1661] = 8'hcc;
 buffer[1662] = 8'h78;
 buffer[1663] = 8'h00;
 buffer[1664] = 8'h00;
 buffer[1665] = 8'h00;
 buffer[1666] = 8'he0;
 buffer[1667] = 8'h60;
 buffer[1668] = 8'h60;
 buffer[1669] = 8'h6c;
 buffer[1670] = 8'h76;
 buffer[1671] = 8'h66;
 buffer[1672] = 8'h66;
 buffer[1673] = 8'h66;
 buffer[1674] = 8'h66;
 buffer[1675] = 8'he6;
 buffer[1676] = 8'h00;
 buffer[1677] = 8'h00;
 buffer[1678] = 8'h00;
 buffer[1679] = 8'h00;
 buffer[1680] = 8'h00;
 buffer[1681] = 8'h00;
 buffer[1682] = 8'h18;
 buffer[1683] = 8'h18;
 buffer[1684] = 8'h00;
 buffer[1685] = 8'h38;
 buffer[1686] = 8'h18;
 buffer[1687] = 8'h18;
 buffer[1688] = 8'h18;
 buffer[1689] = 8'h18;
 buffer[1690] = 8'h18;
 buffer[1691] = 8'h3c;
 buffer[1692] = 8'h00;
 buffer[1693] = 8'h00;
 buffer[1694] = 8'h00;
 buffer[1695] = 8'h00;
 buffer[1696] = 8'h00;
 buffer[1697] = 8'h00;
 buffer[1698] = 8'h06;
 buffer[1699] = 8'h06;
 buffer[1700] = 8'h00;
 buffer[1701] = 8'h0e;
 buffer[1702] = 8'h06;
 buffer[1703] = 8'h06;
 buffer[1704] = 8'h06;
 buffer[1705] = 8'h06;
 buffer[1706] = 8'h06;
 buffer[1707] = 8'h06;
 buffer[1708] = 8'h66;
 buffer[1709] = 8'h66;
 buffer[1710] = 8'h3c;
 buffer[1711] = 8'h00;
 buffer[1712] = 8'h00;
 buffer[1713] = 8'h00;
 buffer[1714] = 8'he0;
 buffer[1715] = 8'h60;
 buffer[1716] = 8'h60;
 buffer[1717] = 8'h66;
 buffer[1718] = 8'h6c;
 buffer[1719] = 8'h78;
 buffer[1720] = 8'h78;
 buffer[1721] = 8'h6c;
 buffer[1722] = 8'h66;
 buffer[1723] = 8'he6;
 buffer[1724] = 8'h00;
 buffer[1725] = 8'h00;
 buffer[1726] = 8'h00;
 buffer[1727] = 8'h00;
 buffer[1728] = 8'h00;
 buffer[1729] = 8'h00;
 buffer[1730] = 8'h38;
 buffer[1731] = 8'h18;
 buffer[1732] = 8'h18;
 buffer[1733] = 8'h18;
 buffer[1734] = 8'h18;
 buffer[1735] = 8'h18;
 buffer[1736] = 8'h18;
 buffer[1737] = 8'h18;
 buffer[1738] = 8'h18;
 buffer[1739] = 8'h3c;
 buffer[1740] = 8'h00;
 buffer[1741] = 8'h00;
 buffer[1742] = 8'h00;
 buffer[1743] = 8'h00;
 buffer[1744] = 8'h00;
 buffer[1745] = 8'h00;
 buffer[1746] = 8'h00;
 buffer[1747] = 8'h00;
 buffer[1748] = 8'h00;
 buffer[1749] = 8'hec;
 buffer[1750] = 8'hfe;
 buffer[1751] = 8'hd6;
 buffer[1752] = 8'hd6;
 buffer[1753] = 8'hd6;
 buffer[1754] = 8'hd6;
 buffer[1755] = 8'hc6;
 buffer[1756] = 8'h00;
 buffer[1757] = 8'h00;
 buffer[1758] = 8'h00;
 buffer[1759] = 8'h00;
 buffer[1760] = 8'h00;
 buffer[1761] = 8'h00;
 buffer[1762] = 8'h00;
 buffer[1763] = 8'h00;
 buffer[1764] = 8'h00;
 buffer[1765] = 8'hdc;
 buffer[1766] = 8'h66;
 buffer[1767] = 8'h66;
 buffer[1768] = 8'h66;
 buffer[1769] = 8'h66;
 buffer[1770] = 8'h66;
 buffer[1771] = 8'h66;
 buffer[1772] = 8'h00;
 buffer[1773] = 8'h00;
 buffer[1774] = 8'h00;
 buffer[1775] = 8'h00;
 buffer[1776] = 8'h00;
 buffer[1777] = 8'h00;
 buffer[1778] = 8'h00;
 buffer[1779] = 8'h00;
 buffer[1780] = 8'h00;
 buffer[1781] = 8'h7c;
 buffer[1782] = 8'hc6;
 buffer[1783] = 8'hc6;
 buffer[1784] = 8'hc6;
 buffer[1785] = 8'hc6;
 buffer[1786] = 8'hc6;
 buffer[1787] = 8'h7c;
 buffer[1788] = 8'h00;
 buffer[1789] = 8'h00;
 buffer[1790] = 8'h00;
 buffer[1791] = 8'h00;
 buffer[1792] = 8'h00;
 buffer[1793] = 8'h00;
 buffer[1794] = 8'h00;
 buffer[1795] = 8'h00;
 buffer[1796] = 8'h00;
 buffer[1797] = 8'hdc;
 buffer[1798] = 8'h66;
 buffer[1799] = 8'h66;
 buffer[1800] = 8'h66;
 buffer[1801] = 8'h66;
 buffer[1802] = 8'h66;
 buffer[1803] = 8'h7c;
 buffer[1804] = 8'h60;
 buffer[1805] = 8'h60;
 buffer[1806] = 8'hf0;
 buffer[1807] = 8'h00;
 buffer[1808] = 8'h00;
 buffer[1809] = 8'h00;
 buffer[1810] = 8'h00;
 buffer[1811] = 8'h00;
 buffer[1812] = 8'h00;
 buffer[1813] = 8'h76;
 buffer[1814] = 8'hcc;
 buffer[1815] = 8'hcc;
 buffer[1816] = 8'hcc;
 buffer[1817] = 8'hcc;
 buffer[1818] = 8'hcc;
 buffer[1819] = 8'h7c;
 buffer[1820] = 8'h0c;
 buffer[1821] = 8'h0c;
 buffer[1822] = 8'h1e;
 buffer[1823] = 8'h00;
 buffer[1824] = 8'h00;
 buffer[1825] = 8'h00;
 buffer[1826] = 8'h00;
 buffer[1827] = 8'h00;
 buffer[1828] = 8'h00;
 buffer[1829] = 8'hdc;
 buffer[1830] = 8'h76;
 buffer[1831] = 8'h66;
 buffer[1832] = 8'h60;
 buffer[1833] = 8'h60;
 buffer[1834] = 8'h60;
 buffer[1835] = 8'hf0;
 buffer[1836] = 8'h00;
 buffer[1837] = 8'h00;
 buffer[1838] = 8'h00;
 buffer[1839] = 8'h00;
 buffer[1840] = 8'h00;
 buffer[1841] = 8'h00;
 buffer[1842] = 8'h00;
 buffer[1843] = 8'h00;
 buffer[1844] = 8'h00;
 buffer[1845] = 8'h7c;
 buffer[1846] = 8'hc6;
 buffer[1847] = 8'h60;
 buffer[1848] = 8'h38;
 buffer[1849] = 8'h0c;
 buffer[1850] = 8'hc6;
 buffer[1851] = 8'h7c;
 buffer[1852] = 8'h00;
 buffer[1853] = 8'h00;
 buffer[1854] = 8'h00;
 buffer[1855] = 8'h00;
 buffer[1856] = 8'h00;
 buffer[1857] = 8'h00;
 buffer[1858] = 8'h10;
 buffer[1859] = 8'h30;
 buffer[1860] = 8'h30;
 buffer[1861] = 8'hfc;
 buffer[1862] = 8'h30;
 buffer[1863] = 8'h30;
 buffer[1864] = 8'h30;
 buffer[1865] = 8'h30;
 buffer[1866] = 8'h36;
 buffer[1867] = 8'h1c;
 buffer[1868] = 8'h00;
 buffer[1869] = 8'h00;
 buffer[1870] = 8'h00;
 buffer[1871] = 8'h00;
 buffer[1872] = 8'h00;
 buffer[1873] = 8'h00;
 buffer[1874] = 8'h00;
 buffer[1875] = 8'h00;
 buffer[1876] = 8'h00;
 buffer[1877] = 8'hcc;
 buffer[1878] = 8'hcc;
 buffer[1879] = 8'hcc;
 buffer[1880] = 8'hcc;
 buffer[1881] = 8'hcc;
 buffer[1882] = 8'hcc;
 buffer[1883] = 8'h76;
 buffer[1884] = 8'h00;
 buffer[1885] = 8'h00;
 buffer[1886] = 8'h00;
 buffer[1887] = 8'h00;
 buffer[1888] = 8'h00;
 buffer[1889] = 8'h00;
 buffer[1890] = 8'h00;
 buffer[1891] = 8'h00;
 buffer[1892] = 8'h00;
 buffer[1893] = 8'h66;
 buffer[1894] = 8'h66;
 buffer[1895] = 8'h66;
 buffer[1896] = 8'h66;
 buffer[1897] = 8'h66;
 buffer[1898] = 8'h3c;
 buffer[1899] = 8'h18;
 buffer[1900] = 8'h00;
 buffer[1901] = 8'h00;
 buffer[1902] = 8'h00;
 buffer[1903] = 8'h00;
 buffer[1904] = 8'h00;
 buffer[1905] = 8'h00;
 buffer[1906] = 8'h00;
 buffer[1907] = 8'h00;
 buffer[1908] = 8'h00;
 buffer[1909] = 8'hc6;
 buffer[1910] = 8'hc6;
 buffer[1911] = 8'hd6;
 buffer[1912] = 8'hd6;
 buffer[1913] = 8'hd6;
 buffer[1914] = 8'hfe;
 buffer[1915] = 8'h6c;
 buffer[1916] = 8'h00;
 buffer[1917] = 8'h00;
 buffer[1918] = 8'h00;
 buffer[1919] = 8'h00;
 buffer[1920] = 8'h00;
 buffer[1921] = 8'h00;
 buffer[1922] = 8'h00;
 buffer[1923] = 8'h00;
 buffer[1924] = 8'h00;
 buffer[1925] = 8'hc6;
 buffer[1926] = 8'h6c;
 buffer[1927] = 8'h38;
 buffer[1928] = 8'h38;
 buffer[1929] = 8'h38;
 buffer[1930] = 8'h6c;
 buffer[1931] = 8'hc6;
 buffer[1932] = 8'h00;
 buffer[1933] = 8'h00;
 buffer[1934] = 8'h00;
 buffer[1935] = 8'h00;
 buffer[1936] = 8'h00;
 buffer[1937] = 8'h00;
 buffer[1938] = 8'h00;
 buffer[1939] = 8'h00;
 buffer[1940] = 8'h00;
 buffer[1941] = 8'hc6;
 buffer[1942] = 8'hc6;
 buffer[1943] = 8'hc6;
 buffer[1944] = 8'hc6;
 buffer[1945] = 8'hc6;
 buffer[1946] = 8'hc6;
 buffer[1947] = 8'h7e;
 buffer[1948] = 8'h06;
 buffer[1949] = 8'h0c;
 buffer[1950] = 8'hf8;
 buffer[1951] = 8'h00;
 buffer[1952] = 8'h00;
 buffer[1953] = 8'h00;
 buffer[1954] = 8'h00;
 buffer[1955] = 8'h00;
 buffer[1956] = 8'h00;
 buffer[1957] = 8'hfe;
 buffer[1958] = 8'hcc;
 buffer[1959] = 8'h18;
 buffer[1960] = 8'h30;
 buffer[1961] = 8'h60;
 buffer[1962] = 8'hc6;
 buffer[1963] = 8'hfe;
 buffer[1964] = 8'h00;
 buffer[1965] = 8'h00;
 buffer[1966] = 8'h00;
 buffer[1967] = 8'h00;
 buffer[1968] = 8'h00;
 buffer[1969] = 8'h00;
 buffer[1970] = 8'h0e;
 buffer[1971] = 8'h18;
 buffer[1972] = 8'h18;
 buffer[1973] = 8'h18;
 buffer[1974] = 8'h70;
 buffer[1975] = 8'h18;
 buffer[1976] = 8'h18;
 buffer[1977] = 8'h18;
 buffer[1978] = 8'h18;
 buffer[1979] = 8'h0e;
 buffer[1980] = 8'h00;
 buffer[1981] = 8'h00;
 buffer[1982] = 8'h00;
 buffer[1983] = 8'h00;
 buffer[1984] = 8'h00;
 buffer[1985] = 8'h00;
 buffer[1986] = 8'h18;
 buffer[1987] = 8'h18;
 buffer[1988] = 8'h18;
 buffer[1989] = 8'h18;
 buffer[1990] = 8'h00;
 buffer[1991] = 8'h18;
 buffer[1992] = 8'h18;
 buffer[1993] = 8'h18;
 buffer[1994] = 8'h18;
 buffer[1995] = 8'h18;
 buffer[1996] = 8'h00;
 buffer[1997] = 8'h00;
 buffer[1998] = 8'h00;
 buffer[1999] = 8'h00;
 buffer[2000] = 8'h00;
 buffer[2001] = 8'h00;
 buffer[2002] = 8'h70;
 buffer[2003] = 8'h18;
 buffer[2004] = 8'h18;
 buffer[2005] = 8'h18;
 buffer[2006] = 8'h0e;
 buffer[2007] = 8'h18;
 buffer[2008] = 8'h18;
 buffer[2009] = 8'h18;
 buffer[2010] = 8'h18;
 buffer[2011] = 8'h70;
 buffer[2012] = 8'h00;
 buffer[2013] = 8'h00;
 buffer[2014] = 8'h00;
 buffer[2015] = 8'h00;
 buffer[2016] = 8'h00;
 buffer[2017] = 8'h00;
 buffer[2018] = 8'h76;
 buffer[2019] = 8'hdc;
 buffer[2020] = 8'h00;
 buffer[2021] = 8'h00;
 buffer[2022] = 8'h00;
 buffer[2023] = 8'h00;
 buffer[2024] = 8'h00;
 buffer[2025] = 8'h00;
 buffer[2026] = 8'h00;
 buffer[2027] = 8'h00;
 buffer[2028] = 8'h00;
 buffer[2029] = 8'h00;
 buffer[2030] = 8'h00;
 buffer[2031] = 8'h00;
 buffer[2032] = 8'h00;
 buffer[2033] = 8'h00;
 buffer[2034] = 8'h00;
 buffer[2035] = 8'h00;
 buffer[2036] = 8'h10;
 buffer[2037] = 8'h38;
 buffer[2038] = 8'h6c;
 buffer[2039] = 8'hc6;
 buffer[2040] = 8'hc6;
 buffer[2041] = 8'hc6;
 buffer[2042] = 8'hfe;
 buffer[2043] = 8'h00;
 buffer[2044] = 8'h00;
 buffer[2045] = 8'h00;
 buffer[2046] = 8'h00;
 buffer[2047] = 8'h00;
 buffer[2048] = 8'h00;
 buffer[2049] = 8'h00;
 buffer[2050] = 8'h3c;
 buffer[2051] = 8'h66;
 buffer[2052] = 8'hc2;
 buffer[2053] = 8'hc0;
 buffer[2054] = 8'hc0;
 buffer[2055] = 8'hc0;
 buffer[2056] = 8'hc2;
 buffer[2057] = 8'h66;
 buffer[2058] = 8'h3c;
 buffer[2059] = 8'h0c;
 buffer[2060] = 8'h06;
 buffer[2061] = 8'h7c;
 buffer[2062] = 8'h00;
 buffer[2063] = 8'h00;
 buffer[2064] = 8'h00;
 buffer[2065] = 8'h00;
 buffer[2066] = 8'hcc;
 buffer[2067] = 8'h00;
 buffer[2068] = 8'h00;
 buffer[2069] = 8'hcc;
 buffer[2070] = 8'hcc;
 buffer[2071] = 8'hcc;
 buffer[2072] = 8'hcc;
 buffer[2073] = 8'hcc;
 buffer[2074] = 8'hcc;
 buffer[2075] = 8'h76;
 buffer[2076] = 8'h00;
 buffer[2077] = 8'h00;
 buffer[2078] = 8'h00;
 buffer[2079] = 8'h00;
 buffer[2080] = 8'h00;
 buffer[2081] = 8'h0c;
 buffer[2082] = 8'h18;
 buffer[2083] = 8'h30;
 buffer[2084] = 8'h00;
 buffer[2085] = 8'h7c;
 buffer[2086] = 8'hc6;
 buffer[2087] = 8'hfe;
 buffer[2088] = 8'hc0;
 buffer[2089] = 8'hc0;
 buffer[2090] = 8'hc6;
 buffer[2091] = 8'h7c;
 buffer[2092] = 8'h00;
 buffer[2093] = 8'h00;
 buffer[2094] = 8'h00;
 buffer[2095] = 8'h00;
 buffer[2096] = 8'h00;
 buffer[2097] = 8'h10;
 buffer[2098] = 8'h38;
 buffer[2099] = 8'h6c;
 buffer[2100] = 8'h00;
 buffer[2101] = 8'h78;
 buffer[2102] = 8'h0c;
 buffer[2103] = 8'h7c;
 buffer[2104] = 8'hcc;
 buffer[2105] = 8'hcc;
 buffer[2106] = 8'hcc;
 buffer[2107] = 8'h76;
 buffer[2108] = 8'h00;
 buffer[2109] = 8'h00;
 buffer[2110] = 8'h00;
 buffer[2111] = 8'h00;
 buffer[2112] = 8'h00;
 buffer[2113] = 8'h00;
 buffer[2114] = 8'hcc;
 buffer[2115] = 8'h00;
 buffer[2116] = 8'h00;
 buffer[2117] = 8'h78;
 buffer[2118] = 8'h0c;
 buffer[2119] = 8'h7c;
 buffer[2120] = 8'hcc;
 buffer[2121] = 8'hcc;
 buffer[2122] = 8'hcc;
 buffer[2123] = 8'h76;
 buffer[2124] = 8'h00;
 buffer[2125] = 8'h00;
 buffer[2126] = 8'h00;
 buffer[2127] = 8'h00;
 buffer[2128] = 8'h00;
 buffer[2129] = 8'h60;
 buffer[2130] = 8'h30;
 buffer[2131] = 8'h18;
 buffer[2132] = 8'h00;
 buffer[2133] = 8'h78;
 buffer[2134] = 8'h0c;
 buffer[2135] = 8'h7c;
 buffer[2136] = 8'hcc;
 buffer[2137] = 8'hcc;
 buffer[2138] = 8'hcc;
 buffer[2139] = 8'h76;
 buffer[2140] = 8'h00;
 buffer[2141] = 8'h00;
 buffer[2142] = 8'h00;
 buffer[2143] = 8'h00;
 buffer[2144] = 8'h00;
 buffer[2145] = 8'h38;
 buffer[2146] = 8'h6c;
 buffer[2147] = 8'h38;
 buffer[2148] = 8'h00;
 buffer[2149] = 8'h78;
 buffer[2150] = 8'h0c;
 buffer[2151] = 8'h7c;
 buffer[2152] = 8'hcc;
 buffer[2153] = 8'hcc;
 buffer[2154] = 8'hcc;
 buffer[2155] = 8'h76;
 buffer[2156] = 8'h00;
 buffer[2157] = 8'h00;
 buffer[2158] = 8'h00;
 buffer[2159] = 8'h00;
 buffer[2160] = 8'h00;
 buffer[2161] = 8'h00;
 buffer[2162] = 8'h00;
 buffer[2163] = 8'h00;
 buffer[2164] = 8'h3c;
 buffer[2165] = 8'h66;
 buffer[2166] = 8'h60;
 buffer[2167] = 8'h60;
 buffer[2168] = 8'h66;
 buffer[2169] = 8'h3c;
 buffer[2170] = 8'h0c;
 buffer[2171] = 8'h06;
 buffer[2172] = 8'h3c;
 buffer[2173] = 8'h00;
 buffer[2174] = 8'h00;
 buffer[2175] = 8'h00;
 buffer[2176] = 8'h00;
 buffer[2177] = 8'h10;
 buffer[2178] = 8'h38;
 buffer[2179] = 8'h6c;
 buffer[2180] = 8'h00;
 buffer[2181] = 8'h7c;
 buffer[2182] = 8'hc6;
 buffer[2183] = 8'hfe;
 buffer[2184] = 8'hc0;
 buffer[2185] = 8'hc0;
 buffer[2186] = 8'hc6;
 buffer[2187] = 8'h7c;
 buffer[2188] = 8'h00;
 buffer[2189] = 8'h00;
 buffer[2190] = 8'h00;
 buffer[2191] = 8'h00;
 buffer[2192] = 8'h00;
 buffer[2193] = 8'h00;
 buffer[2194] = 8'hc6;
 buffer[2195] = 8'h00;
 buffer[2196] = 8'h00;
 buffer[2197] = 8'h7c;
 buffer[2198] = 8'hc6;
 buffer[2199] = 8'hfe;
 buffer[2200] = 8'hc0;
 buffer[2201] = 8'hc0;
 buffer[2202] = 8'hc6;
 buffer[2203] = 8'h7c;
 buffer[2204] = 8'h00;
 buffer[2205] = 8'h00;
 buffer[2206] = 8'h00;
 buffer[2207] = 8'h00;
 buffer[2208] = 8'h00;
 buffer[2209] = 8'h60;
 buffer[2210] = 8'h30;
 buffer[2211] = 8'h18;
 buffer[2212] = 8'h00;
 buffer[2213] = 8'h7c;
 buffer[2214] = 8'hc6;
 buffer[2215] = 8'hfe;
 buffer[2216] = 8'hc0;
 buffer[2217] = 8'hc0;
 buffer[2218] = 8'hc6;
 buffer[2219] = 8'h7c;
 buffer[2220] = 8'h00;
 buffer[2221] = 8'h00;
 buffer[2222] = 8'h00;
 buffer[2223] = 8'h00;
 buffer[2224] = 8'h00;
 buffer[2225] = 8'h00;
 buffer[2226] = 8'h66;
 buffer[2227] = 8'h00;
 buffer[2228] = 8'h00;
 buffer[2229] = 8'h38;
 buffer[2230] = 8'h18;
 buffer[2231] = 8'h18;
 buffer[2232] = 8'h18;
 buffer[2233] = 8'h18;
 buffer[2234] = 8'h18;
 buffer[2235] = 8'h3c;
 buffer[2236] = 8'h00;
 buffer[2237] = 8'h00;
 buffer[2238] = 8'h00;
 buffer[2239] = 8'h00;
 buffer[2240] = 8'h00;
 buffer[2241] = 8'h18;
 buffer[2242] = 8'h3c;
 buffer[2243] = 8'h66;
 buffer[2244] = 8'h00;
 buffer[2245] = 8'h38;
 buffer[2246] = 8'h18;
 buffer[2247] = 8'h18;
 buffer[2248] = 8'h18;
 buffer[2249] = 8'h18;
 buffer[2250] = 8'h18;
 buffer[2251] = 8'h3c;
 buffer[2252] = 8'h00;
 buffer[2253] = 8'h00;
 buffer[2254] = 8'h00;
 buffer[2255] = 8'h00;
 buffer[2256] = 8'h00;
 buffer[2257] = 8'h60;
 buffer[2258] = 8'h30;
 buffer[2259] = 8'h18;
 buffer[2260] = 8'h00;
 buffer[2261] = 8'h38;
 buffer[2262] = 8'h18;
 buffer[2263] = 8'h18;
 buffer[2264] = 8'h18;
 buffer[2265] = 8'h18;
 buffer[2266] = 8'h18;
 buffer[2267] = 8'h3c;
 buffer[2268] = 8'h00;
 buffer[2269] = 8'h00;
 buffer[2270] = 8'h00;
 buffer[2271] = 8'h00;
 buffer[2272] = 8'h00;
 buffer[2273] = 8'hc6;
 buffer[2274] = 8'h00;
 buffer[2275] = 8'h10;
 buffer[2276] = 8'h38;
 buffer[2277] = 8'h6c;
 buffer[2278] = 8'hc6;
 buffer[2279] = 8'hc6;
 buffer[2280] = 8'hfe;
 buffer[2281] = 8'hc6;
 buffer[2282] = 8'hc6;
 buffer[2283] = 8'hc6;
 buffer[2284] = 8'h00;
 buffer[2285] = 8'h00;
 buffer[2286] = 8'h00;
 buffer[2287] = 8'h00;
 buffer[2288] = 8'h38;
 buffer[2289] = 8'h6c;
 buffer[2290] = 8'h38;
 buffer[2291] = 8'h00;
 buffer[2292] = 8'h38;
 buffer[2293] = 8'h6c;
 buffer[2294] = 8'hc6;
 buffer[2295] = 8'hc6;
 buffer[2296] = 8'hfe;
 buffer[2297] = 8'hc6;
 buffer[2298] = 8'hc6;
 buffer[2299] = 8'hc6;
 buffer[2300] = 8'h00;
 buffer[2301] = 8'h00;
 buffer[2302] = 8'h00;
 buffer[2303] = 8'h00;
 buffer[2304] = 8'h18;
 buffer[2305] = 8'h30;
 buffer[2306] = 8'h60;
 buffer[2307] = 8'h00;
 buffer[2308] = 8'hfe;
 buffer[2309] = 8'h66;
 buffer[2310] = 8'h60;
 buffer[2311] = 8'h7c;
 buffer[2312] = 8'h60;
 buffer[2313] = 8'h60;
 buffer[2314] = 8'h66;
 buffer[2315] = 8'hfe;
 buffer[2316] = 8'h00;
 buffer[2317] = 8'h00;
 buffer[2318] = 8'h00;
 buffer[2319] = 8'h00;
 buffer[2320] = 8'h00;
 buffer[2321] = 8'h00;
 buffer[2322] = 8'h00;
 buffer[2323] = 8'h00;
 buffer[2324] = 8'h00;
 buffer[2325] = 8'hcc;
 buffer[2326] = 8'h76;
 buffer[2327] = 8'h36;
 buffer[2328] = 8'h7e;
 buffer[2329] = 8'hd8;
 buffer[2330] = 8'hd8;
 buffer[2331] = 8'h6e;
 buffer[2332] = 8'h00;
 buffer[2333] = 8'h00;
 buffer[2334] = 8'h00;
 buffer[2335] = 8'h00;
 buffer[2336] = 8'h00;
 buffer[2337] = 8'h00;
 buffer[2338] = 8'h3e;
 buffer[2339] = 8'h6c;
 buffer[2340] = 8'hcc;
 buffer[2341] = 8'hcc;
 buffer[2342] = 8'hfe;
 buffer[2343] = 8'hcc;
 buffer[2344] = 8'hcc;
 buffer[2345] = 8'hcc;
 buffer[2346] = 8'hcc;
 buffer[2347] = 8'hce;
 buffer[2348] = 8'h00;
 buffer[2349] = 8'h00;
 buffer[2350] = 8'h00;
 buffer[2351] = 8'h00;
 buffer[2352] = 8'h00;
 buffer[2353] = 8'h10;
 buffer[2354] = 8'h38;
 buffer[2355] = 8'h6c;
 buffer[2356] = 8'h00;
 buffer[2357] = 8'h7c;
 buffer[2358] = 8'hc6;
 buffer[2359] = 8'hc6;
 buffer[2360] = 8'hc6;
 buffer[2361] = 8'hc6;
 buffer[2362] = 8'hc6;
 buffer[2363] = 8'h7c;
 buffer[2364] = 8'h00;
 buffer[2365] = 8'h00;
 buffer[2366] = 8'h00;
 buffer[2367] = 8'h00;
 buffer[2368] = 8'h00;
 buffer[2369] = 8'h00;
 buffer[2370] = 8'hc6;
 buffer[2371] = 8'h00;
 buffer[2372] = 8'h00;
 buffer[2373] = 8'h7c;
 buffer[2374] = 8'hc6;
 buffer[2375] = 8'hc6;
 buffer[2376] = 8'hc6;
 buffer[2377] = 8'hc6;
 buffer[2378] = 8'hc6;
 buffer[2379] = 8'h7c;
 buffer[2380] = 8'h00;
 buffer[2381] = 8'h00;
 buffer[2382] = 8'h00;
 buffer[2383] = 8'h00;
 buffer[2384] = 8'h00;
 buffer[2385] = 8'h60;
 buffer[2386] = 8'h30;
 buffer[2387] = 8'h18;
 buffer[2388] = 8'h00;
 buffer[2389] = 8'h7c;
 buffer[2390] = 8'hc6;
 buffer[2391] = 8'hc6;
 buffer[2392] = 8'hc6;
 buffer[2393] = 8'hc6;
 buffer[2394] = 8'hc6;
 buffer[2395] = 8'h7c;
 buffer[2396] = 8'h00;
 buffer[2397] = 8'h00;
 buffer[2398] = 8'h00;
 buffer[2399] = 8'h00;
 buffer[2400] = 8'h00;
 buffer[2401] = 8'h30;
 buffer[2402] = 8'h78;
 buffer[2403] = 8'hcc;
 buffer[2404] = 8'h00;
 buffer[2405] = 8'hcc;
 buffer[2406] = 8'hcc;
 buffer[2407] = 8'hcc;
 buffer[2408] = 8'hcc;
 buffer[2409] = 8'hcc;
 buffer[2410] = 8'hcc;
 buffer[2411] = 8'h76;
 buffer[2412] = 8'h00;
 buffer[2413] = 8'h00;
 buffer[2414] = 8'h00;
 buffer[2415] = 8'h00;
 buffer[2416] = 8'h00;
 buffer[2417] = 8'h60;
 buffer[2418] = 8'h30;
 buffer[2419] = 8'h18;
 buffer[2420] = 8'h00;
 buffer[2421] = 8'hcc;
 buffer[2422] = 8'hcc;
 buffer[2423] = 8'hcc;
 buffer[2424] = 8'hcc;
 buffer[2425] = 8'hcc;
 buffer[2426] = 8'hcc;
 buffer[2427] = 8'h76;
 buffer[2428] = 8'h00;
 buffer[2429] = 8'h00;
 buffer[2430] = 8'h00;
 buffer[2431] = 8'h00;
 buffer[2432] = 8'h00;
 buffer[2433] = 8'h00;
 buffer[2434] = 8'hc6;
 buffer[2435] = 8'h00;
 buffer[2436] = 8'h00;
 buffer[2437] = 8'hc6;
 buffer[2438] = 8'hc6;
 buffer[2439] = 8'hc6;
 buffer[2440] = 8'hc6;
 buffer[2441] = 8'hc6;
 buffer[2442] = 8'hc6;
 buffer[2443] = 8'h7e;
 buffer[2444] = 8'h06;
 buffer[2445] = 8'h0c;
 buffer[2446] = 8'h78;
 buffer[2447] = 8'h00;
 buffer[2448] = 8'h00;
 buffer[2449] = 8'hc6;
 buffer[2450] = 8'h00;
 buffer[2451] = 8'h7c;
 buffer[2452] = 8'hc6;
 buffer[2453] = 8'hc6;
 buffer[2454] = 8'hc6;
 buffer[2455] = 8'hc6;
 buffer[2456] = 8'hc6;
 buffer[2457] = 8'hc6;
 buffer[2458] = 8'hc6;
 buffer[2459] = 8'h7c;
 buffer[2460] = 8'h00;
 buffer[2461] = 8'h00;
 buffer[2462] = 8'h00;
 buffer[2463] = 8'h00;
 buffer[2464] = 8'h00;
 buffer[2465] = 8'hc6;
 buffer[2466] = 8'h00;
 buffer[2467] = 8'hc6;
 buffer[2468] = 8'hc6;
 buffer[2469] = 8'hc6;
 buffer[2470] = 8'hc6;
 buffer[2471] = 8'hc6;
 buffer[2472] = 8'hc6;
 buffer[2473] = 8'hc6;
 buffer[2474] = 8'hc6;
 buffer[2475] = 8'h7c;
 buffer[2476] = 8'h00;
 buffer[2477] = 8'h00;
 buffer[2478] = 8'h00;
 buffer[2479] = 8'h00;
 buffer[2480] = 8'h00;
 buffer[2481] = 8'h18;
 buffer[2482] = 8'h18;
 buffer[2483] = 8'h3c;
 buffer[2484] = 8'h66;
 buffer[2485] = 8'h60;
 buffer[2486] = 8'h60;
 buffer[2487] = 8'h60;
 buffer[2488] = 8'h66;
 buffer[2489] = 8'h3c;
 buffer[2490] = 8'h18;
 buffer[2491] = 8'h18;
 buffer[2492] = 8'h00;
 buffer[2493] = 8'h00;
 buffer[2494] = 8'h00;
 buffer[2495] = 8'h00;
 buffer[2496] = 8'h00;
 buffer[2497] = 8'h38;
 buffer[2498] = 8'h6c;
 buffer[2499] = 8'h64;
 buffer[2500] = 8'h60;
 buffer[2501] = 8'hf0;
 buffer[2502] = 8'h60;
 buffer[2503] = 8'h60;
 buffer[2504] = 8'h60;
 buffer[2505] = 8'h60;
 buffer[2506] = 8'he6;
 buffer[2507] = 8'hfc;
 buffer[2508] = 8'h00;
 buffer[2509] = 8'h00;
 buffer[2510] = 8'h00;
 buffer[2511] = 8'h00;
 buffer[2512] = 8'h00;
 buffer[2513] = 8'h00;
 buffer[2514] = 8'h66;
 buffer[2515] = 8'h66;
 buffer[2516] = 8'h3c;
 buffer[2517] = 8'h18;
 buffer[2518] = 8'h7e;
 buffer[2519] = 8'h18;
 buffer[2520] = 8'h7e;
 buffer[2521] = 8'h18;
 buffer[2522] = 8'h18;
 buffer[2523] = 8'h18;
 buffer[2524] = 8'h00;
 buffer[2525] = 8'h00;
 buffer[2526] = 8'h00;
 buffer[2527] = 8'h00;
 buffer[2528] = 8'h00;
 buffer[2529] = 8'hf8;
 buffer[2530] = 8'hcc;
 buffer[2531] = 8'hcc;
 buffer[2532] = 8'hf8;
 buffer[2533] = 8'hc4;
 buffer[2534] = 8'hcc;
 buffer[2535] = 8'hde;
 buffer[2536] = 8'hcc;
 buffer[2537] = 8'hcc;
 buffer[2538] = 8'hcc;
 buffer[2539] = 8'hc6;
 buffer[2540] = 8'h00;
 buffer[2541] = 8'h00;
 buffer[2542] = 8'h00;
 buffer[2543] = 8'h00;
 buffer[2544] = 8'h00;
 buffer[2545] = 8'h0e;
 buffer[2546] = 8'h1b;
 buffer[2547] = 8'h18;
 buffer[2548] = 8'h18;
 buffer[2549] = 8'h18;
 buffer[2550] = 8'h7e;
 buffer[2551] = 8'h18;
 buffer[2552] = 8'h18;
 buffer[2553] = 8'h18;
 buffer[2554] = 8'h18;
 buffer[2555] = 8'h18;
 buffer[2556] = 8'hd8;
 buffer[2557] = 8'h70;
 buffer[2558] = 8'h00;
 buffer[2559] = 8'h00;
 buffer[2560] = 8'h00;
 buffer[2561] = 8'h18;
 buffer[2562] = 8'h30;
 buffer[2563] = 8'h60;
 buffer[2564] = 8'h00;
 buffer[2565] = 8'h78;
 buffer[2566] = 8'h0c;
 buffer[2567] = 8'h7c;
 buffer[2568] = 8'hcc;
 buffer[2569] = 8'hcc;
 buffer[2570] = 8'hcc;
 buffer[2571] = 8'h76;
 buffer[2572] = 8'h00;
 buffer[2573] = 8'h00;
 buffer[2574] = 8'h00;
 buffer[2575] = 8'h00;
 buffer[2576] = 8'h00;
 buffer[2577] = 8'h0c;
 buffer[2578] = 8'h18;
 buffer[2579] = 8'h30;
 buffer[2580] = 8'h00;
 buffer[2581] = 8'h38;
 buffer[2582] = 8'h18;
 buffer[2583] = 8'h18;
 buffer[2584] = 8'h18;
 buffer[2585] = 8'h18;
 buffer[2586] = 8'h18;
 buffer[2587] = 8'h3c;
 buffer[2588] = 8'h00;
 buffer[2589] = 8'h00;
 buffer[2590] = 8'h00;
 buffer[2591] = 8'h00;
 buffer[2592] = 8'h00;
 buffer[2593] = 8'h18;
 buffer[2594] = 8'h30;
 buffer[2595] = 8'h60;
 buffer[2596] = 8'h00;
 buffer[2597] = 8'h7c;
 buffer[2598] = 8'hc6;
 buffer[2599] = 8'hc6;
 buffer[2600] = 8'hc6;
 buffer[2601] = 8'hc6;
 buffer[2602] = 8'hc6;
 buffer[2603] = 8'h7c;
 buffer[2604] = 8'h00;
 buffer[2605] = 8'h00;
 buffer[2606] = 8'h00;
 buffer[2607] = 8'h00;
 buffer[2608] = 8'h00;
 buffer[2609] = 8'h18;
 buffer[2610] = 8'h30;
 buffer[2611] = 8'h60;
 buffer[2612] = 8'h00;
 buffer[2613] = 8'hcc;
 buffer[2614] = 8'hcc;
 buffer[2615] = 8'hcc;
 buffer[2616] = 8'hcc;
 buffer[2617] = 8'hcc;
 buffer[2618] = 8'hcc;
 buffer[2619] = 8'h76;
 buffer[2620] = 8'h00;
 buffer[2621] = 8'h00;
 buffer[2622] = 8'h00;
 buffer[2623] = 8'h00;
 buffer[2624] = 8'h00;
 buffer[2625] = 8'h00;
 buffer[2626] = 8'h76;
 buffer[2627] = 8'hdc;
 buffer[2628] = 8'h00;
 buffer[2629] = 8'hdc;
 buffer[2630] = 8'h66;
 buffer[2631] = 8'h66;
 buffer[2632] = 8'h66;
 buffer[2633] = 8'h66;
 buffer[2634] = 8'h66;
 buffer[2635] = 8'h66;
 buffer[2636] = 8'h00;
 buffer[2637] = 8'h00;
 buffer[2638] = 8'h00;
 buffer[2639] = 8'h00;
 buffer[2640] = 8'h76;
 buffer[2641] = 8'hdc;
 buffer[2642] = 8'h00;
 buffer[2643] = 8'hc6;
 buffer[2644] = 8'he6;
 buffer[2645] = 8'hf6;
 buffer[2646] = 8'hfe;
 buffer[2647] = 8'hde;
 buffer[2648] = 8'hce;
 buffer[2649] = 8'hc6;
 buffer[2650] = 8'hc6;
 buffer[2651] = 8'hc6;
 buffer[2652] = 8'h00;
 buffer[2653] = 8'h00;
 buffer[2654] = 8'h00;
 buffer[2655] = 8'h00;
 buffer[2656] = 8'h00;
 buffer[2657] = 8'h3c;
 buffer[2658] = 8'h6c;
 buffer[2659] = 8'h6c;
 buffer[2660] = 8'h3e;
 buffer[2661] = 8'h00;
 buffer[2662] = 8'h7e;
 buffer[2663] = 8'h00;
 buffer[2664] = 8'h00;
 buffer[2665] = 8'h00;
 buffer[2666] = 8'h00;
 buffer[2667] = 8'h00;
 buffer[2668] = 8'h00;
 buffer[2669] = 8'h00;
 buffer[2670] = 8'h00;
 buffer[2671] = 8'h00;
 buffer[2672] = 8'h00;
 buffer[2673] = 8'h38;
 buffer[2674] = 8'h6c;
 buffer[2675] = 8'h6c;
 buffer[2676] = 8'h38;
 buffer[2677] = 8'h00;
 buffer[2678] = 8'h7c;
 buffer[2679] = 8'h00;
 buffer[2680] = 8'h00;
 buffer[2681] = 8'h00;
 buffer[2682] = 8'h00;
 buffer[2683] = 8'h00;
 buffer[2684] = 8'h00;
 buffer[2685] = 8'h00;
 buffer[2686] = 8'h00;
 buffer[2687] = 8'h00;
 buffer[2688] = 8'h00;
 buffer[2689] = 8'h00;
 buffer[2690] = 8'h30;
 buffer[2691] = 8'h30;
 buffer[2692] = 8'h00;
 buffer[2693] = 8'h30;
 buffer[2694] = 8'h30;
 buffer[2695] = 8'h60;
 buffer[2696] = 8'hc0;
 buffer[2697] = 8'hc6;
 buffer[2698] = 8'hc6;
 buffer[2699] = 8'h7c;
 buffer[2700] = 8'h00;
 buffer[2701] = 8'h00;
 buffer[2702] = 8'h00;
 buffer[2703] = 8'h00;
 buffer[2704] = 8'h00;
 buffer[2705] = 8'h00;
 buffer[2706] = 8'h00;
 buffer[2707] = 8'h00;
 buffer[2708] = 8'h00;
 buffer[2709] = 8'h00;
 buffer[2710] = 8'hfe;
 buffer[2711] = 8'hc0;
 buffer[2712] = 8'hc0;
 buffer[2713] = 8'hc0;
 buffer[2714] = 8'hc0;
 buffer[2715] = 8'h00;
 buffer[2716] = 8'h00;
 buffer[2717] = 8'h00;
 buffer[2718] = 8'h00;
 buffer[2719] = 8'h00;
 buffer[2720] = 8'h00;
 buffer[2721] = 8'h00;
 buffer[2722] = 8'h00;
 buffer[2723] = 8'h00;
 buffer[2724] = 8'h00;
 buffer[2725] = 8'h00;
 buffer[2726] = 8'hfe;
 buffer[2727] = 8'h06;
 buffer[2728] = 8'h06;
 buffer[2729] = 8'h06;
 buffer[2730] = 8'h06;
 buffer[2731] = 8'h00;
 buffer[2732] = 8'h00;
 buffer[2733] = 8'h00;
 buffer[2734] = 8'h00;
 buffer[2735] = 8'h00;
 buffer[2736] = 8'h00;
 buffer[2737] = 8'hc0;
 buffer[2738] = 8'hc0;
 buffer[2739] = 8'hc2;
 buffer[2740] = 8'hc6;
 buffer[2741] = 8'hcc;
 buffer[2742] = 8'h18;
 buffer[2743] = 8'h30;
 buffer[2744] = 8'h60;
 buffer[2745] = 8'hdc;
 buffer[2746] = 8'h86;
 buffer[2747] = 8'h0c;
 buffer[2748] = 8'h18;
 buffer[2749] = 8'h3e;
 buffer[2750] = 8'h00;
 buffer[2751] = 8'h00;
 buffer[2752] = 8'h00;
 buffer[2753] = 8'hc0;
 buffer[2754] = 8'hc0;
 buffer[2755] = 8'hc2;
 buffer[2756] = 8'hc6;
 buffer[2757] = 8'hcc;
 buffer[2758] = 8'h18;
 buffer[2759] = 8'h30;
 buffer[2760] = 8'h66;
 buffer[2761] = 8'hce;
 buffer[2762] = 8'h9e;
 buffer[2763] = 8'h3e;
 buffer[2764] = 8'h06;
 buffer[2765] = 8'h06;
 buffer[2766] = 8'h00;
 buffer[2767] = 8'h00;
 buffer[2768] = 8'h00;
 buffer[2769] = 8'h00;
 buffer[2770] = 8'h18;
 buffer[2771] = 8'h18;
 buffer[2772] = 8'h00;
 buffer[2773] = 8'h18;
 buffer[2774] = 8'h18;
 buffer[2775] = 8'h18;
 buffer[2776] = 8'h3c;
 buffer[2777] = 8'h3c;
 buffer[2778] = 8'h3c;
 buffer[2779] = 8'h18;
 buffer[2780] = 8'h00;
 buffer[2781] = 8'h00;
 buffer[2782] = 8'h00;
 buffer[2783] = 8'h00;
 buffer[2784] = 8'h00;
 buffer[2785] = 8'h00;
 buffer[2786] = 8'h00;
 buffer[2787] = 8'h00;
 buffer[2788] = 8'h00;
 buffer[2789] = 8'h36;
 buffer[2790] = 8'h6c;
 buffer[2791] = 8'hd8;
 buffer[2792] = 8'h6c;
 buffer[2793] = 8'h36;
 buffer[2794] = 8'h00;
 buffer[2795] = 8'h00;
 buffer[2796] = 8'h00;
 buffer[2797] = 8'h00;
 buffer[2798] = 8'h00;
 buffer[2799] = 8'h00;
 buffer[2800] = 8'h00;
 buffer[2801] = 8'h00;
 buffer[2802] = 8'h00;
 buffer[2803] = 8'h00;
 buffer[2804] = 8'h00;
 buffer[2805] = 8'hd8;
 buffer[2806] = 8'h6c;
 buffer[2807] = 8'h36;
 buffer[2808] = 8'h6c;
 buffer[2809] = 8'hd8;
 buffer[2810] = 8'h00;
 buffer[2811] = 8'h00;
 buffer[2812] = 8'h00;
 buffer[2813] = 8'h00;
 buffer[2814] = 8'h00;
 buffer[2815] = 8'h00;
 buffer[2816] = 8'h11;
 buffer[2817] = 8'h44;
 buffer[2818] = 8'h11;
 buffer[2819] = 8'h44;
 buffer[2820] = 8'h11;
 buffer[2821] = 8'h44;
 buffer[2822] = 8'h11;
 buffer[2823] = 8'h44;
 buffer[2824] = 8'h11;
 buffer[2825] = 8'h44;
 buffer[2826] = 8'h11;
 buffer[2827] = 8'h44;
 buffer[2828] = 8'h11;
 buffer[2829] = 8'h44;
 buffer[2830] = 8'h11;
 buffer[2831] = 8'h44;
 buffer[2832] = 8'h55;
 buffer[2833] = 8'haa;
 buffer[2834] = 8'h55;
 buffer[2835] = 8'haa;
 buffer[2836] = 8'h55;
 buffer[2837] = 8'haa;
 buffer[2838] = 8'h55;
 buffer[2839] = 8'haa;
 buffer[2840] = 8'h55;
 buffer[2841] = 8'haa;
 buffer[2842] = 8'h55;
 buffer[2843] = 8'haa;
 buffer[2844] = 8'h55;
 buffer[2845] = 8'haa;
 buffer[2846] = 8'h55;
 buffer[2847] = 8'haa;
 buffer[2848] = 8'hdd;
 buffer[2849] = 8'h77;
 buffer[2850] = 8'hdd;
 buffer[2851] = 8'h77;
 buffer[2852] = 8'hdd;
 buffer[2853] = 8'h77;
 buffer[2854] = 8'hdd;
 buffer[2855] = 8'h77;
 buffer[2856] = 8'hdd;
 buffer[2857] = 8'h77;
 buffer[2858] = 8'hdd;
 buffer[2859] = 8'h77;
 buffer[2860] = 8'hdd;
 buffer[2861] = 8'h77;
 buffer[2862] = 8'hdd;
 buffer[2863] = 8'h77;
 buffer[2864] = 8'h18;
 buffer[2865] = 8'h18;
 buffer[2866] = 8'h18;
 buffer[2867] = 8'h18;
 buffer[2868] = 8'h18;
 buffer[2869] = 8'h18;
 buffer[2870] = 8'h18;
 buffer[2871] = 8'h18;
 buffer[2872] = 8'h18;
 buffer[2873] = 8'h18;
 buffer[2874] = 8'h18;
 buffer[2875] = 8'h18;
 buffer[2876] = 8'h18;
 buffer[2877] = 8'h18;
 buffer[2878] = 8'h18;
 buffer[2879] = 8'h18;
 buffer[2880] = 8'h18;
 buffer[2881] = 8'h18;
 buffer[2882] = 8'h18;
 buffer[2883] = 8'h18;
 buffer[2884] = 8'h18;
 buffer[2885] = 8'h18;
 buffer[2886] = 8'h18;
 buffer[2887] = 8'hf8;
 buffer[2888] = 8'h18;
 buffer[2889] = 8'h18;
 buffer[2890] = 8'h18;
 buffer[2891] = 8'h18;
 buffer[2892] = 8'h18;
 buffer[2893] = 8'h18;
 buffer[2894] = 8'h18;
 buffer[2895] = 8'h18;
 buffer[2896] = 8'h18;
 buffer[2897] = 8'h18;
 buffer[2898] = 8'h18;
 buffer[2899] = 8'h18;
 buffer[2900] = 8'h18;
 buffer[2901] = 8'hf8;
 buffer[2902] = 8'h18;
 buffer[2903] = 8'hf8;
 buffer[2904] = 8'h18;
 buffer[2905] = 8'h18;
 buffer[2906] = 8'h18;
 buffer[2907] = 8'h18;
 buffer[2908] = 8'h18;
 buffer[2909] = 8'h18;
 buffer[2910] = 8'h18;
 buffer[2911] = 8'h18;
 buffer[2912] = 8'h36;
 buffer[2913] = 8'h36;
 buffer[2914] = 8'h36;
 buffer[2915] = 8'h36;
 buffer[2916] = 8'h36;
 buffer[2917] = 8'h36;
 buffer[2918] = 8'h36;
 buffer[2919] = 8'hf6;
 buffer[2920] = 8'h36;
 buffer[2921] = 8'h36;
 buffer[2922] = 8'h36;
 buffer[2923] = 8'h36;
 buffer[2924] = 8'h36;
 buffer[2925] = 8'h36;
 buffer[2926] = 8'h36;
 buffer[2927] = 8'h36;
 buffer[2928] = 8'h00;
 buffer[2929] = 8'h00;
 buffer[2930] = 8'h00;
 buffer[2931] = 8'h00;
 buffer[2932] = 8'h00;
 buffer[2933] = 8'h00;
 buffer[2934] = 8'h00;
 buffer[2935] = 8'hfe;
 buffer[2936] = 8'h36;
 buffer[2937] = 8'h36;
 buffer[2938] = 8'h36;
 buffer[2939] = 8'h36;
 buffer[2940] = 8'h36;
 buffer[2941] = 8'h36;
 buffer[2942] = 8'h36;
 buffer[2943] = 8'h36;
 buffer[2944] = 8'h00;
 buffer[2945] = 8'h00;
 buffer[2946] = 8'h00;
 buffer[2947] = 8'h00;
 buffer[2948] = 8'h00;
 buffer[2949] = 8'hf8;
 buffer[2950] = 8'h18;
 buffer[2951] = 8'hf8;
 buffer[2952] = 8'h18;
 buffer[2953] = 8'h18;
 buffer[2954] = 8'h18;
 buffer[2955] = 8'h18;
 buffer[2956] = 8'h18;
 buffer[2957] = 8'h18;
 buffer[2958] = 8'h18;
 buffer[2959] = 8'h18;
 buffer[2960] = 8'h36;
 buffer[2961] = 8'h36;
 buffer[2962] = 8'h36;
 buffer[2963] = 8'h36;
 buffer[2964] = 8'h36;
 buffer[2965] = 8'hf6;
 buffer[2966] = 8'h06;
 buffer[2967] = 8'hf6;
 buffer[2968] = 8'h36;
 buffer[2969] = 8'h36;
 buffer[2970] = 8'h36;
 buffer[2971] = 8'h36;
 buffer[2972] = 8'h36;
 buffer[2973] = 8'h36;
 buffer[2974] = 8'h36;
 buffer[2975] = 8'h36;
 buffer[2976] = 8'h36;
 buffer[2977] = 8'h36;
 buffer[2978] = 8'h36;
 buffer[2979] = 8'h36;
 buffer[2980] = 8'h36;
 buffer[2981] = 8'h36;
 buffer[2982] = 8'h36;
 buffer[2983] = 8'h36;
 buffer[2984] = 8'h36;
 buffer[2985] = 8'h36;
 buffer[2986] = 8'h36;
 buffer[2987] = 8'h36;
 buffer[2988] = 8'h36;
 buffer[2989] = 8'h36;
 buffer[2990] = 8'h36;
 buffer[2991] = 8'h36;
 buffer[2992] = 8'h00;
 buffer[2993] = 8'h00;
 buffer[2994] = 8'h00;
 buffer[2995] = 8'h00;
 buffer[2996] = 8'h00;
 buffer[2997] = 8'hfe;
 buffer[2998] = 8'h06;
 buffer[2999] = 8'hf6;
 buffer[3000] = 8'h36;
 buffer[3001] = 8'h36;
 buffer[3002] = 8'h36;
 buffer[3003] = 8'h36;
 buffer[3004] = 8'h36;
 buffer[3005] = 8'h36;
 buffer[3006] = 8'h36;
 buffer[3007] = 8'h36;
 buffer[3008] = 8'h36;
 buffer[3009] = 8'h36;
 buffer[3010] = 8'h36;
 buffer[3011] = 8'h36;
 buffer[3012] = 8'h36;
 buffer[3013] = 8'hf6;
 buffer[3014] = 8'h06;
 buffer[3015] = 8'hfe;
 buffer[3016] = 8'h00;
 buffer[3017] = 8'h00;
 buffer[3018] = 8'h00;
 buffer[3019] = 8'h00;
 buffer[3020] = 8'h00;
 buffer[3021] = 8'h00;
 buffer[3022] = 8'h00;
 buffer[3023] = 8'h00;
 buffer[3024] = 8'h36;
 buffer[3025] = 8'h36;
 buffer[3026] = 8'h36;
 buffer[3027] = 8'h36;
 buffer[3028] = 8'h36;
 buffer[3029] = 8'h36;
 buffer[3030] = 8'h36;
 buffer[3031] = 8'hfe;
 buffer[3032] = 8'h00;
 buffer[3033] = 8'h00;
 buffer[3034] = 8'h00;
 buffer[3035] = 8'h00;
 buffer[3036] = 8'h00;
 buffer[3037] = 8'h00;
 buffer[3038] = 8'h00;
 buffer[3039] = 8'h00;
 buffer[3040] = 8'h18;
 buffer[3041] = 8'h18;
 buffer[3042] = 8'h18;
 buffer[3043] = 8'h18;
 buffer[3044] = 8'h18;
 buffer[3045] = 8'hf8;
 buffer[3046] = 8'h18;
 buffer[3047] = 8'hf8;
 buffer[3048] = 8'h00;
 buffer[3049] = 8'h00;
 buffer[3050] = 8'h00;
 buffer[3051] = 8'h00;
 buffer[3052] = 8'h00;
 buffer[3053] = 8'h00;
 buffer[3054] = 8'h00;
 buffer[3055] = 8'h00;
 buffer[3056] = 8'h00;
 buffer[3057] = 8'h00;
 buffer[3058] = 8'h00;
 buffer[3059] = 8'h00;
 buffer[3060] = 8'h00;
 buffer[3061] = 8'h00;
 buffer[3062] = 8'h00;
 buffer[3063] = 8'hf8;
 buffer[3064] = 8'h18;
 buffer[3065] = 8'h18;
 buffer[3066] = 8'h18;
 buffer[3067] = 8'h18;
 buffer[3068] = 8'h18;
 buffer[3069] = 8'h18;
 buffer[3070] = 8'h18;
 buffer[3071] = 8'h18;
 buffer[3072] = 8'h18;
 buffer[3073] = 8'h18;
 buffer[3074] = 8'h18;
 buffer[3075] = 8'h18;
 buffer[3076] = 8'h18;
 buffer[3077] = 8'h18;
 buffer[3078] = 8'h18;
 buffer[3079] = 8'h1f;
 buffer[3080] = 8'h00;
 buffer[3081] = 8'h00;
 buffer[3082] = 8'h00;
 buffer[3083] = 8'h00;
 buffer[3084] = 8'h00;
 buffer[3085] = 8'h00;
 buffer[3086] = 8'h00;
 buffer[3087] = 8'h00;
 buffer[3088] = 8'h18;
 buffer[3089] = 8'h18;
 buffer[3090] = 8'h18;
 buffer[3091] = 8'h18;
 buffer[3092] = 8'h18;
 buffer[3093] = 8'h18;
 buffer[3094] = 8'h18;
 buffer[3095] = 8'hff;
 buffer[3096] = 8'h00;
 buffer[3097] = 8'h00;
 buffer[3098] = 8'h00;
 buffer[3099] = 8'h00;
 buffer[3100] = 8'h00;
 buffer[3101] = 8'h00;
 buffer[3102] = 8'h00;
 buffer[3103] = 8'h00;
 buffer[3104] = 8'h00;
 buffer[3105] = 8'h00;
 buffer[3106] = 8'h00;
 buffer[3107] = 8'h00;
 buffer[3108] = 8'h00;
 buffer[3109] = 8'h00;
 buffer[3110] = 8'h00;
 buffer[3111] = 8'hff;
 buffer[3112] = 8'h18;
 buffer[3113] = 8'h18;
 buffer[3114] = 8'h18;
 buffer[3115] = 8'h18;
 buffer[3116] = 8'h18;
 buffer[3117] = 8'h18;
 buffer[3118] = 8'h18;
 buffer[3119] = 8'h18;
 buffer[3120] = 8'h18;
 buffer[3121] = 8'h18;
 buffer[3122] = 8'h18;
 buffer[3123] = 8'h18;
 buffer[3124] = 8'h18;
 buffer[3125] = 8'h18;
 buffer[3126] = 8'h18;
 buffer[3127] = 8'h1f;
 buffer[3128] = 8'h18;
 buffer[3129] = 8'h18;
 buffer[3130] = 8'h18;
 buffer[3131] = 8'h18;
 buffer[3132] = 8'h18;
 buffer[3133] = 8'h18;
 buffer[3134] = 8'h18;
 buffer[3135] = 8'h18;
 buffer[3136] = 8'h00;
 buffer[3137] = 8'h00;
 buffer[3138] = 8'h00;
 buffer[3139] = 8'h00;
 buffer[3140] = 8'h00;
 buffer[3141] = 8'h00;
 buffer[3142] = 8'h00;
 buffer[3143] = 8'hff;
 buffer[3144] = 8'h00;
 buffer[3145] = 8'h00;
 buffer[3146] = 8'h00;
 buffer[3147] = 8'h00;
 buffer[3148] = 8'h00;
 buffer[3149] = 8'h00;
 buffer[3150] = 8'h00;
 buffer[3151] = 8'h00;
 buffer[3152] = 8'h18;
 buffer[3153] = 8'h18;
 buffer[3154] = 8'h18;
 buffer[3155] = 8'h18;
 buffer[3156] = 8'h18;
 buffer[3157] = 8'h18;
 buffer[3158] = 8'h18;
 buffer[3159] = 8'hff;
 buffer[3160] = 8'h18;
 buffer[3161] = 8'h18;
 buffer[3162] = 8'h18;
 buffer[3163] = 8'h18;
 buffer[3164] = 8'h18;
 buffer[3165] = 8'h18;
 buffer[3166] = 8'h18;
 buffer[3167] = 8'h18;
 buffer[3168] = 8'h18;
 buffer[3169] = 8'h18;
 buffer[3170] = 8'h18;
 buffer[3171] = 8'h18;
 buffer[3172] = 8'h18;
 buffer[3173] = 8'h1f;
 buffer[3174] = 8'h18;
 buffer[3175] = 8'h1f;
 buffer[3176] = 8'h18;
 buffer[3177] = 8'h18;
 buffer[3178] = 8'h18;
 buffer[3179] = 8'h18;
 buffer[3180] = 8'h18;
 buffer[3181] = 8'h18;
 buffer[3182] = 8'h18;
 buffer[3183] = 8'h18;
 buffer[3184] = 8'h36;
 buffer[3185] = 8'h36;
 buffer[3186] = 8'h36;
 buffer[3187] = 8'h36;
 buffer[3188] = 8'h36;
 buffer[3189] = 8'h36;
 buffer[3190] = 8'h36;
 buffer[3191] = 8'h37;
 buffer[3192] = 8'h36;
 buffer[3193] = 8'h36;
 buffer[3194] = 8'h36;
 buffer[3195] = 8'h36;
 buffer[3196] = 8'h36;
 buffer[3197] = 8'h36;
 buffer[3198] = 8'h36;
 buffer[3199] = 8'h36;
 buffer[3200] = 8'h36;
 buffer[3201] = 8'h36;
 buffer[3202] = 8'h36;
 buffer[3203] = 8'h36;
 buffer[3204] = 8'h36;
 buffer[3205] = 8'h37;
 buffer[3206] = 8'h30;
 buffer[3207] = 8'h3f;
 buffer[3208] = 8'h00;
 buffer[3209] = 8'h00;
 buffer[3210] = 8'h00;
 buffer[3211] = 8'h00;
 buffer[3212] = 8'h00;
 buffer[3213] = 8'h00;
 buffer[3214] = 8'h00;
 buffer[3215] = 8'h00;
 buffer[3216] = 8'h00;
 buffer[3217] = 8'h00;
 buffer[3218] = 8'h00;
 buffer[3219] = 8'h00;
 buffer[3220] = 8'h00;
 buffer[3221] = 8'h3f;
 buffer[3222] = 8'h30;
 buffer[3223] = 8'h37;
 buffer[3224] = 8'h36;
 buffer[3225] = 8'h36;
 buffer[3226] = 8'h36;
 buffer[3227] = 8'h36;
 buffer[3228] = 8'h36;
 buffer[3229] = 8'h36;
 buffer[3230] = 8'h36;
 buffer[3231] = 8'h36;
 buffer[3232] = 8'h36;
 buffer[3233] = 8'h36;
 buffer[3234] = 8'h36;
 buffer[3235] = 8'h36;
 buffer[3236] = 8'h36;
 buffer[3237] = 8'hf7;
 buffer[3238] = 8'h00;
 buffer[3239] = 8'hff;
 buffer[3240] = 8'h00;
 buffer[3241] = 8'h00;
 buffer[3242] = 8'h00;
 buffer[3243] = 8'h00;
 buffer[3244] = 8'h00;
 buffer[3245] = 8'h00;
 buffer[3246] = 8'h00;
 buffer[3247] = 8'h00;
 buffer[3248] = 8'h00;
 buffer[3249] = 8'h00;
 buffer[3250] = 8'h00;
 buffer[3251] = 8'h00;
 buffer[3252] = 8'h00;
 buffer[3253] = 8'hff;
 buffer[3254] = 8'h00;
 buffer[3255] = 8'hf7;
 buffer[3256] = 8'h36;
 buffer[3257] = 8'h36;
 buffer[3258] = 8'h36;
 buffer[3259] = 8'h36;
 buffer[3260] = 8'h36;
 buffer[3261] = 8'h36;
 buffer[3262] = 8'h36;
 buffer[3263] = 8'h36;
 buffer[3264] = 8'h36;
 buffer[3265] = 8'h36;
 buffer[3266] = 8'h36;
 buffer[3267] = 8'h36;
 buffer[3268] = 8'h36;
 buffer[3269] = 8'h37;
 buffer[3270] = 8'h30;
 buffer[3271] = 8'h37;
 buffer[3272] = 8'h36;
 buffer[3273] = 8'h36;
 buffer[3274] = 8'h36;
 buffer[3275] = 8'h36;
 buffer[3276] = 8'h36;
 buffer[3277] = 8'h36;
 buffer[3278] = 8'h36;
 buffer[3279] = 8'h36;
 buffer[3280] = 8'h00;
 buffer[3281] = 8'h00;
 buffer[3282] = 8'h00;
 buffer[3283] = 8'h00;
 buffer[3284] = 8'h00;
 buffer[3285] = 8'hff;
 buffer[3286] = 8'h00;
 buffer[3287] = 8'hff;
 buffer[3288] = 8'h00;
 buffer[3289] = 8'h00;
 buffer[3290] = 8'h00;
 buffer[3291] = 8'h00;
 buffer[3292] = 8'h00;
 buffer[3293] = 8'h00;
 buffer[3294] = 8'h00;
 buffer[3295] = 8'h00;
 buffer[3296] = 8'h36;
 buffer[3297] = 8'h36;
 buffer[3298] = 8'h36;
 buffer[3299] = 8'h36;
 buffer[3300] = 8'h36;
 buffer[3301] = 8'hf7;
 buffer[3302] = 8'h00;
 buffer[3303] = 8'hf7;
 buffer[3304] = 8'h36;
 buffer[3305] = 8'h36;
 buffer[3306] = 8'h36;
 buffer[3307] = 8'h36;
 buffer[3308] = 8'h36;
 buffer[3309] = 8'h36;
 buffer[3310] = 8'h36;
 buffer[3311] = 8'h36;
 buffer[3312] = 8'h18;
 buffer[3313] = 8'h18;
 buffer[3314] = 8'h18;
 buffer[3315] = 8'h18;
 buffer[3316] = 8'h18;
 buffer[3317] = 8'hff;
 buffer[3318] = 8'h00;
 buffer[3319] = 8'hff;
 buffer[3320] = 8'h00;
 buffer[3321] = 8'h00;
 buffer[3322] = 8'h00;
 buffer[3323] = 8'h00;
 buffer[3324] = 8'h00;
 buffer[3325] = 8'h00;
 buffer[3326] = 8'h00;
 buffer[3327] = 8'h00;
 buffer[3328] = 8'h36;
 buffer[3329] = 8'h36;
 buffer[3330] = 8'h36;
 buffer[3331] = 8'h36;
 buffer[3332] = 8'h36;
 buffer[3333] = 8'h36;
 buffer[3334] = 8'h36;
 buffer[3335] = 8'hff;
 buffer[3336] = 8'h00;
 buffer[3337] = 8'h00;
 buffer[3338] = 8'h00;
 buffer[3339] = 8'h00;
 buffer[3340] = 8'h00;
 buffer[3341] = 8'h00;
 buffer[3342] = 8'h00;
 buffer[3343] = 8'h00;
 buffer[3344] = 8'h00;
 buffer[3345] = 8'h00;
 buffer[3346] = 8'h00;
 buffer[3347] = 8'h00;
 buffer[3348] = 8'h00;
 buffer[3349] = 8'hff;
 buffer[3350] = 8'h00;
 buffer[3351] = 8'hff;
 buffer[3352] = 8'h18;
 buffer[3353] = 8'h18;
 buffer[3354] = 8'h18;
 buffer[3355] = 8'h18;
 buffer[3356] = 8'h18;
 buffer[3357] = 8'h18;
 buffer[3358] = 8'h18;
 buffer[3359] = 8'h18;
 buffer[3360] = 8'h00;
 buffer[3361] = 8'h00;
 buffer[3362] = 8'h00;
 buffer[3363] = 8'h00;
 buffer[3364] = 8'h00;
 buffer[3365] = 8'h00;
 buffer[3366] = 8'h00;
 buffer[3367] = 8'hff;
 buffer[3368] = 8'h36;
 buffer[3369] = 8'h36;
 buffer[3370] = 8'h36;
 buffer[3371] = 8'h36;
 buffer[3372] = 8'h36;
 buffer[3373] = 8'h36;
 buffer[3374] = 8'h36;
 buffer[3375] = 8'h36;
 buffer[3376] = 8'h36;
 buffer[3377] = 8'h36;
 buffer[3378] = 8'h36;
 buffer[3379] = 8'h36;
 buffer[3380] = 8'h36;
 buffer[3381] = 8'h36;
 buffer[3382] = 8'h36;
 buffer[3383] = 8'h3f;
 buffer[3384] = 8'h00;
 buffer[3385] = 8'h00;
 buffer[3386] = 8'h00;
 buffer[3387] = 8'h00;
 buffer[3388] = 8'h00;
 buffer[3389] = 8'h00;
 buffer[3390] = 8'h00;
 buffer[3391] = 8'h00;
 buffer[3392] = 8'h18;
 buffer[3393] = 8'h18;
 buffer[3394] = 8'h18;
 buffer[3395] = 8'h18;
 buffer[3396] = 8'h18;
 buffer[3397] = 8'h1f;
 buffer[3398] = 8'h18;
 buffer[3399] = 8'h1f;
 buffer[3400] = 8'h00;
 buffer[3401] = 8'h00;
 buffer[3402] = 8'h00;
 buffer[3403] = 8'h00;
 buffer[3404] = 8'h00;
 buffer[3405] = 8'h00;
 buffer[3406] = 8'h00;
 buffer[3407] = 8'h00;
 buffer[3408] = 8'h00;
 buffer[3409] = 8'h00;
 buffer[3410] = 8'h00;
 buffer[3411] = 8'h00;
 buffer[3412] = 8'h00;
 buffer[3413] = 8'h1f;
 buffer[3414] = 8'h18;
 buffer[3415] = 8'h1f;
 buffer[3416] = 8'h18;
 buffer[3417] = 8'h18;
 buffer[3418] = 8'h18;
 buffer[3419] = 8'h18;
 buffer[3420] = 8'h18;
 buffer[3421] = 8'h18;
 buffer[3422] = 8'h18;
 buffer[3423] = 8'h18;
 buffer[3424] = 8'h00;
 buffer[3425] = 8'h00;
 buffer[3426] = 8'h00;
 buffer[3427] = 8'h00;
 buffer[3428] = 8'h00;
 buffer[3429] = 8'h00;
 buffer[3430] = 8'h00;
 buffer[3431] = 8'h3f;
 buffer[3432] = 8'h36;
 buffer[3433] = 8'h36;
 buffer[3434] = 8'h36;
 buffer[3435] = 8'h36;
 buffer[3436] = 8'h36;
 buffer[3437] = 8'h36;
 buffer[3438] = 8'h36;
 buffer[3439] = 8'h36;
 buffer[3440] = 8'h36;
 buffer[3441] = 8'h36;
 buffer[3442] = 8'h36;
 buffer[3443] = 8'h36;
 buffer[3444] = 8'h36;
 buffer[3445] = 8'h36;
 buffer[3446] = 8'h36;
 buffer[3447] = 8'hff;
 buffer[3448] = 8'h36;
 buffer[3449] = 8'h36;
 buffer[3450] = 8'h36;
 buffer[3451] = 8'h36;
 buffer[3452] = 8'h36;
 buffer[3453] = 8'h36;
 buffer[3454] = 8'h36;
 buffer[3455] = 8'h36;
 buffer[3456] = 8'h18;
 buffer[3457] = 8'h18;
 buffer[3458] = 8'h18;
 buffer[3459] = 8'h18;
 buffer[3460] = 8'h18;
 buffer[3461] = 8'hff;
 buffer[3462] = 8'h18;
 buffer[3463] = 8'hff;
 buffer[3464] = 8'h18;
 buffer[3465] = 8'h18;
 buffer[3466] = 8'h18;
 buffer[3467] = 8'h18;
 buffer[3468] = 8'h18;
 buffer[3469] = 8'h18;
 buffer[3470] = 8'h18;
 buffer[3471] = 8'h18;
 buffer[3472] = 8'h18;
 buffer[3473] = 8'h18;
 buffer[3474] = 8'h18;
 buffer[3475] = 8'h18;
 buffer[3476] = 8'h18;
 buffer[3477] = 8'h18;
 buffer[3478] = 8'h18;
 buffer[3479] = 8'hf8;
 buffer[3480] = 8'h00;
 buffer[3481] = 8'h00;
 buffer[3482] = 8'h00;
 buffer[3483] = 8'h00;
 buffer[3484] = 8'h00;
 buffer[3485] = 8'h00;
 buffer[3486] = 8'h00;
 buffer[3487] = 8'h00;
 buffer[3488] = 8'h00;
 buffer[3489] = 8'h00;
 buffer[3490] = 8'h00;
 buffer[3491] = 8'h00;
 buffer[3492] = 8'h00;
 buffer[3493] = 8'h00;
 buffer[3494] = 8'h00;
 buffer[3495] = 8'h1f;
 buffer[3496] = 8'h18;
 buffer[3497] = 8'h18;
 buffer[3498] = 8'h18;
 buffer[3499] = 8'h18;
 buffer[3500] = 8'h18;
 buffer[3501] = 8'h18;
 buffer[3502] = 8'h18;
 buffer[3503] = 8'h18;
 buffer[3504] = 8'hff;
 buffer[3505] = 8'hff;
 buffer[3506] = 8'hff;
 buffer[3507] = 8'hff;
 buffer[3508] = 8'hff;
 buffer[3509] = 8'hff;
 buffer[3510] = 8'hff;
 buffer[3511] = 8'hff;
 buffer[3512] = 8'hff;
 buffer[3513] = 8'hff;
 buffer[3514] = 8'hff;
 buffer[3515] = 8'hff;
 buffer[3516] = 8'hff;
 buffer[3517] = 8'hff;
 buffer[3518] = 8'hff;
 buffer[3519] = 8'hff;
 buffer[3520] = 8'h00;
 buffer[3521] = 8'h00;
 buffer[3522] = 8'h00;
 buffer[3523] = 8'h00;
 buffer[3524] = 8'h00;
 buffer[3525] = 8'h00;
 buffer[3526] = 8'h00;
 buffer[3527] = 8'hff;
 buffer[3528] = 8'hff;
 buffer[3529] = 8'hff;
 buffer[3530] = 8'hff;
 buffer[3531] = 8'hff;
 buffer[3532] = 8'hff;
 buffer[3533] = 8'hff;
 buffer[3534] = 8'hff;
 buffer[3535] = 8'hff;
 buffer[3536] = 8'hf0;
 buffer[3537] = 8'hf0;
 buffer[3538] = 8'hf0;
 buffer[3539] = 8'hf0;
 buffer[3540] = 8'hf0;
 buffer[3541] = 8'hf0;
 buffer[3542] = 8'hf0;
 buffer[3543] = 8'hf0;
 buffer[3544] = 8'hf0;
 buffer[3545] = 8'hf0;
 buffer[3546] = 8'hf0;
 buffer[3547] = 8'hf0;
 buffer[3548] = 8'hf0;
 buffer[3549] = 8'hf0;
 buffer[3550] = 8'hf0;
 buffer[3551] = 8'hf0;
 buffer[3552] = 8'h0f;
 buffer[3553] = 8'h0f;
 buffer[3554] = 8'h0f;
 buffer[3555] = 8'h0f;
 buffer[3556] = 8'h0f;
 buffer[3557] = 8'h0f;
 buffer[3558] = 8'h0f;
 buffer[3559] = 8'h0f;
 buffer[3560] = 8'h0f;
 buffer[3561] = 8'h0f;
 buffer[3562] = 8'h0f;
 buffer[3563] = 8'h0f;
 buffer[3564] = 8'h0f;
 buffer[3565] = 8'h0f;
 buffer[3566] = 8'h0f;
 buffer[3567] = 8'h0f;
 buffer[3568] = 8'hff;
 buffer[3569] = 8'hff;
 buffer[3570] = 8'hff;
 buffer[3571] = 8'hff;
 buffer[3572] = 8'hff;
 buffer[3573] = 8'hff;
 buffer[3574] = 8'hff;
 buffer[3575] = 8'h00;
 buffer[3576] = 8'h00;
 buffer[3577] = 8'h00;
 buffer[3578] = 8'h00;
 buffer[3579] = 8'h00;
 buffer[3580] = 8'h00;
 buffer[3581] = 8'h00;
 buffer[3582] = 8'h00;
 buffer[3583] = 8'h00;
 buffer[3584] = 8'h00;
 buffer[3585] = 8'h00;
 buffer[3586] = 8'h00;
 buffer[3587] = 8'h00;
 buffer[3588] = 8'h00;
 buffer[3589] = 8'h76;
 buffer[3590] = 8'hdc;
 buffer[3591] = 8'hd8;
 buffer[3592] = 8'hd8;
 buffer[3593] = 8'hd8;
 buffer[3594] = 8'hdc;
 buffer[3595] = 8'h76;
 buffer[3596] = 8'h00;
 buffer[3597] = 8'h00;
 buffer[3598] = 8'h00;
 buffer[3599] = 8'h00;
 buffer[3600] = 8'h00;
 buffer[3601] = 8'h00;
 buffer[3602] = 8'h78;
 buffer[3603] = 8'hcc;
 buffer[3604] = 8'hcc;
 buffer[3605] = 8'hcc;
 buffer[3606] = 8'hd8;
 buffer[3607] = 8'hcc;
 buffer[3608] = 8'hc6;
 buffer[3609] = 8'hc6;
 buffer[3610] = 8'hc6;
 buffer[3611] = 8'hcc;
 buffer[3612] = 8'h00;
 buffer[3613] = 8'h00;
 buffer[3614] = 8'h00;
 buffer[3615] = 8'h00;
 buffer[3616] = 8'h00;
 buffer[3617] = 8'h00;
 buffer[3618] = 8'hfe;
 buffer[3619] = 8'hc6;
 buffer[3620] = 8'hc6;
 buffer[3621] = 8'hc0;
 buffer[3622] = 8'hc0;
 buffer[3623] = 8'hc0;
 buffer[3624] = 8'hc0;
 buffer[3625] = 8'hc0;
 buffer[3626] = 8'hc0;
 buffer[3627] = 8'hc0;
 buffer[3628] = 8'h00;
 buffer[3629] = 8'h00;
 buffer[3630] = 8'h00;
 buffer[3631] = 8'h00;
 buffer[3632] = 8'h00;
 buffer[3633] = 8'h00;
 buffer[3634] = 8'h00;
 buffer[3635] = 8'h00;
 buffer[3636] = 8'hfe;
 buffer[3637] = 8'h6c;
 buffer[3638] = 8'h6c;
 buffer[3639] = 8'h6c;
 buffer[3640] = 8'h6c;
 buffer[3641] = 8'h6c;
 buffer[3642] = 8'h6c;
 buffer[3643] = 8'h6c;
 buffer[3644] = 8'h00;
 buffer[3645] = 8'h00;
 buffer[3646] = 8'h00;
 buffer[3647] = 8'h00;
 buffer[3648] = 8'h00;
 buffer[3649] = 8'h00;
 buffer[3650] = 8'h00;
 buffer[3651] = 8'hfe;
 buffer[3652] = 8'hc6;
 buffer[3653] = 8'h60;
 buffer[3654] = 8'h30;
 buffer[3655] = 8'h18;
 buffer[3656] = 8'h30;
 buffer[3657] = 8'h60;
 buffer[3658] = 8'hc6;
 buffer[3659] = 8'hfe;
 buffer[3660] = 8'h00;
 buffer[3661] = 8'h00;
 buffer[3662] = 8'h00;
 buffer[3663] = 8'h00;
 buffer[3664] = 8'h00;
 buffer[3665] = 8'h00;
 buffer[3666] = 8'h00;
 buffer[3667] = 8'h00;
 buffer[3668] = 8'h00;
 buffer[3669] = 8'h7e;
 buffer[3670] = 8'hd8;
 buffer[3671] = 8'hd8;
 buffer[3672] = 8'hd8;
 buffer[3673] = 8'hd8;
 buffer[3674] = 8'hd8;
 buffer[3675] = 8'h70;
 buffer[3676] = 8'h00;
 buffer[3677] = 8'h00;
 buffer[3678] = 8'h00;
 buffer[3679] = 8'h00;
 buffer[3680] = 8'h00;
 buffer[3681] = 8'h00;
 buffer[3682] = 8'h00;
 buffer[3683] = 8'h00;
 buffer[3684] = 8'h66;
 buffer[3685] = 8'h66;
 buffer[3686] = 8'h66;
 buffer[3687] = 8'h66;
 buffer[3688] = 8'h66;
 buffer[3689] = 8'h7c;
 buffer[3690] = 8'h60;
 buffer[3691] = 8'h60;
 buffer[3692] = 8'hc0;
 buffer[3693] = 8'h00;
 buffer[3694] = 8'h00;
 buffer[3695] = 8'h00;
 buffer[3696] = 8'h00;
 buffer[3697] = 8'h00;
 buffer[3698] = 8'h00;
 buffer[3699] = 8'h00;
 buffer[3700] = 8'h76;
 buffer[3701] = 8'hdc;
 buffer[3702] = 8'h18;
 buffer[3703] = 8'h18;
 buffer[3704] = 8'h18;
 buffer[3705] = 8'h18;
 buffer[3706] = 8'h18;
 buffer[3707] = 8'h18;
 buffer[3708] = 8'h00;
 buffer[3709] = 8'h00;
 buffer[3710] = 8'h00;
 buffer[3711] = 8'h00;
 buffer[3712] = 8'h00;
 buffer[3713] = 8'h00;
 buffer[3714] = 8'h00;
 buffer[3715] = 8'h7e;
 buffer[3716] = 8'h18;
 buffer[3717] = 8'h3c;
 buffer[3718] = 8'h66;
 buffer[3719] = 8'h66;
 buffer[3720] = 8'h66;
 buffer[3721] = 8'h3c;
 buffer[3722] = 8'h18;
 buffer[3723] = 8'h7e;
 buffer[3724] = 8'h00;
 buffer[3725] = 8'h00;
 buffer[3726] = 8'h00;
 buffer[3727] = 8'h00;
 buffer[3728] = 8'h00;
 buffer[3729] = 8'h00;
 buffer[3730] = 8'h00;
 buffer[3731] = 8'h38;
 buffer[3732] = 8'h6c;
 buffer[3733] = 8'hc6;
 buffer[3734] = 8'hc6;
 buffer[3735] = 8'hfe;
 buffer[3736] = 8'hc6;
 buffer[3737] = 8'hc6;
 buffer[3738] = 8'h6c;
 buffer[3739] = 8'h38;
 buffer[3740] = 8'h00;
 buffer[3741] = 8'h00;
 buffer[3742] = 8'h00;
 buffer[3743] = 8'h00;
 buffer[3744] = 8'h00;
 buffer[3745] = 8'h00;
 buffer[3746] = 8'h38;
 buffer[3747] = 8'h6c;
 buffer[3748] = 8'hc6;
 buffer[3749] = 8'hc6;
 buffer[3750] = 8'hc6;
 buffer[3751] = 8'h6c;
 buffer[3752] = 8'h6c;
 buffer[3753] = 8'h6c;
 buffer[3754] = 8'h6c;
 buffer[3755] = 8'hee;
 buffer[3756] = 8'h00;
 buffer[3757] = 8'h00;
 buffer[3758] = 8'h00;
 buffer[3759] = 8'h00;
 buffer[3760] = 8'h00;
 buffer[3761] = 8'h00;
 buffer[3762] = 8'h1e;
 buffer[3763] = 8'h30;
 buffer[3764] = 8'h18;
 buffer[3765] = 8'h0c;
 buffer[3766] = 8'h3e;
 buffer[3767] = 8'h66;
 buffer[3768] = 8'h66;
 buffer[3769] = 8'h66;
 buffer[3770] = 8'h66;
 buffer[3771] = 8'h3c;
 buffer[3772] = 8'h00;
 buffer[3773] = 8'h00;
 buffer[3774] = 8'h00;
 buffer[3775] = 8'h00;
 buffer[3776] = 8'h00;
 buffer[3777] = 8'h00;
 buffer[3778] = 8'h00;
 buffer[3779] = 8'h00;
 buffer[3780] = 8'h00;
 buffer[3781] = 8'h7e;
 buffer[3782] = 8'hdb;
 buffer[3783] = 8'hdb;
 buffer[3784] = 8'hdb;
 buffer[3785] = 8'h7e;
 buffer[3786] = 8'h00;
 buffer[3787] = 8'h00;
 buffer[3788] = 8'h00;
 buffer[3789] = 8'h00;
 buffer[3790] = 8'h00;
 buffer[3791] = 8'h00;
 buffer[3792] = 8'h00;
 buffer[3793] = 8'h00;
 buffer[3794] = 8'h00;
 buffer[3795] = 8'h03;
 buffer[3796] = 8'h06;
 buffer[3797] = 8'h7e;
 buffer[3798] = 8'hdb;
 buffer[3799] = 8'hdb;
 buffer[3800] = 8'hf3;
 buffer[3801] = 8'h7e;
 buffer[3802] = 8'h60;
 buffer[3803] = 8'hc0;
 buffer[3804] = 8'h00;
 buffer[3805] = 8'h00;
 buffer[3806] = 8'h00;
 buffer[3807] = 8'h00;
 buffer[3808] = 8'h00;
 buffer[3809] = 8'h00;
 buffer[3810] = 8'h1c;
 buffer[3811] = 8'h30;
 buffer[3812] = 8'h60;
 buffer[3813] = 8'h60;
 buffer[3814] = 8'h7c;
 buffer[3815] = 8'h60;
 buffer[3816] = 8'h60;
 buffer[3817] = 8'h60;
 buffer[3818] = 8'h30;
 buffer[3819] = 8'h1c;
 buffer[3820] = 8'h00;
 buffer[3821] = 8'h00;
 buffer[3822] = 8'h00;
 buffer[3823] = 8'h00;
 buffer[3824] = 8'h00;
 buffer[3825] = 8'h00;
 buffer[3826] = 8'h00;
 buffer[3827] = 8'h7c;
 buffer[3828] = 8'hc6;
 buffer[3829] = 8'hc6;
 buffer[3830] = 8'hc6;
 buffer[3831] = 8'hc6;
 buffer[3832] = 8'hc6;
 buffer[3833] = 8'hc6;
 buffer[3834] = 8'hc6;
 buffer[3835] = 8'hc6;
 buffer[3836] = 8'h00;
 buffer[3837] = 8'h00;
 buffer[3838] = 8'h00;
 buffer[3839] = 8'h00;
 buffer[3840] = 8'h00;
 buffer[3841] = 8'h00;
 buffer[3842] = 8'h00;
 buffer[3843] = 8'h00;
 buffer[3844] = 8'hfe;
 buffer[3845] = 8'h00;
 buffer[3846] = 8'h00;
 buffer[3847] = 8'hfe;
 buffer[3848] = 8'h00;
 buffer[3849] = 8'h00;
 buffer[3850] = 8'hfe;
 buffer[3851] = 8'h00;
 buffer[3852] = 8'h00;
 buffer[3853] = 8'h00;
 buffer[3854] = 8'h00;
 buffer[3855] = 8'h00;
 buffer[3856] = 8'h00;
 buffer[3857] = 8'h00;
 buffer[3858] = 8'h00;
 buffer[3859] = 8'h00;
 buffer[3860] = 8'h18;
 buffer[3861] = 8'h18;
 buffer[3862] = 8'h7e;
 buffer[3863] = 8'h18;
 buffer[3864] = 8'h18;
 buffer[3865] = 8'h00;
 buffer[3866] = 8'h00;
 buffer[3867] = 8'hff;
 buffer[3868] = 8'h00;
 buffer[3869] = 8'h00;
 buffer[3870] = 8'h00;
 buffer[3871] = 8'h00;
 buffer[3872] = 8'h00;
 buffer[3873] = 8'h00;
 buffer[3874] = 8'h00;
 buffer[3875] = 8'h30;
 buffer[3876] = 8'h18;
 buffer[3877] = 8'h0c;
 buffer[3878] = 8'h06;
 buffer[3879] = 8'h0c;
 buffer[3880] = 8'h18;
 buffer[3881] = 8'h30;
 buffer[3882] = 8'h00;
 buffer[3883] = 8'h7e;
 buffer[3884] = 8'h00;
 buffer[3885] = 8'h00;
 buffer[3886] = 8'h00;
 buffer[3887] = 8'h00;
 buffer[3888] = 8'h00;
 buffer[3889] = 8'h00;
 buffer[3890] = 8'h00;
 buffer[3891] = 8'h0c;
 buffer[3892] = 8'h18;
 buffer[3893] = 8'h30;
 buffer[3894] = 8'h60;
 buffer[3895] = 8'h30;
 buffer[3896] = 8'h18;
 buffer[3897] = 8'h0c;
 buffer[3898] = 8'h00;
 buffer[3899] = 8'h7e;
 buffer[3900] = 8'h00;
 buffer[3901] = 8'h00;
 buffer[3902] = 8'h00;
 buffer[3903] = 8'h00;
 buffer[3904] = 8'h00;
 buffer[3905] = 8'h00;
 buffer[3906] = 8'h0e;
 buffer[3907] = 8'h1b;
 buffer[3908] = 8'h1b;
 buffer[3909] = 8'h18;
 buffer[3910] = 8'h18;
 buffer[3911] = 8'h18;
 buffer[3912] = 8'h18;
 buffer[3913] = 8'h18;
 buffer[3914] = 8'h18;
 buffer[3915] = 8'h18;
 buffer[3916] = 8'h18;
 buffer[3917] = 8'h18;
 buffer[3918] = 8'h18;
 buffer[3919] = 8'h18;
 buffer[3920] = 8'h18;
 buffer[3921] = 8'h18;
 buffer[3922] = 8'h18;
 buffer[3923] = 8'h18;
 buffer[3924] = 8'h18;
 buffer[3925] = 8'h18;
 buffer[3926] = 8'h18;
 buffer[3927] = 8'h18;
 buffer[3928] = 8'hd8;
 buffer[3929] = 8'hd8;
 buffer[3930] = 8'hd8;
 buffer[3931] = 8'h70;
 buffer[3932] = 8'h00;
 buffer[3933] = 8'h00;
 buffer[3934] = 8'h00;
 buffer[3935] = 8'h00;
 buffer[3936] = 8'h00;
 buffer[3937] = 8'h00;
 buffer[3938] = 8'h00;
 buffer[3939] = 8'h00;
 buffer[3940] = 8'h18;
 buffer[3941] = 8'h18;
 buffer[3942] = 8'h00;
 buffer[3943] = 8'h7e;
 buffer[3944] = 8'h00;
 buffer[3945] = 8'h18;
 buffer[3946] = 8'h18;
 buffer[3947] = 8'h00;
 buffer[3948] = 8'h00;
 buffer[3949] = 8'h00;
 buffer[3950] = 8'h00;
 buffer[3951] = 8'h00;
 buffer[3952] = 8'h00;
 buffer[3953] = 8'h00;
 buffer[3954] = 8'h00;
 buffer[3955] = 8'h00;
 buffer[3956] = 8'h00;
 buffer[3957] = 8'h76;
 buffer[3958] = 8'hdc;
 buffer[3959] = 8'h00;
 buffer[3960] = 8'h76;
 buffer[3961] = 8'hdc;
 buffer[3962] = 8'h00;
 buffer[3963] = 8'h00;
 buffer[3964] = 8'h00;
 buffer[3965] = 8'h00;
 buffer[3966] = 8'h00;
 buffer[3967] = 8'h00;
 buffer[3968] = 8'h00;
 buffer[3969] = 8'h38;
 buffer[3970] = 8'h6c;
 buffer[3971] = 8'h6c;
 buffer[3972] = 8'h38;
 buffer[3973] = 8'h00;
 buffer[3974] = 8'h00;
 buffer[3975] = 8'h00;
 buffer[3976] = 8'h00;
 buffer[3977] = 8'h00;
 buffer[3978] = 8'h00;
 buffer[3979] = 8'h00;
 buffer[3980] = 8'h00;
 buffer[3981] = 8'h00;
 buffer[3982] = 8'h00;
 buffer[3983] = 8'h00;
 buffer[3984] = 8'h00;
 buffer[3985] = 8'h00;
 buffer[3986] = 8'h00;
 buffer[3987] = 8'h00;
 buffer[3988] = 8'h00;
 buffer[3989] = 8'h00;
 buffer[3990] = 8'h00;
 buffer[3991] = 8'h18;
 buffer[3992] = 8'h18;
 buffer[3993] = 8'h00;
 buffer[3994] = 8'h00;
 buffer[3995] = 8'h00;
 buffer[3996] = 8'h00;
 buffer[3997] = 8'h00;
 buffer[3998] = 8'h00;
 buffer[3999] = 8'h00;
 buffer[4000] = 8'h00;
 buffer[4001] = 8'h00;
 buffer[4002] = 8'h00;
 buffer[4003] = 8'h00;
 buffer[4004] = 8'h00;
 buffer[4005] = 8'h00;
 buffer[4006] = 8'h00;
 buffer[4007] = 8'h00;
 buffer[4008] = 8'h18;
 buffer[4009] = 8'h00;
 buffer[4010] = 8'h00;
 buffer[4011] = 8'h00;
 buffer[4012] = 8'h00;
 buffer[4013] = 8'h00;
 buffer[4014] = 8'h00;
 buffer[4015] = 8'h00;
 buffer[4016] = 8'h00;
 buffer[4017] = 8'h0f;
 buffer[4018] = 8'h0c;
 buffer[4019] = 8'h0c;
 buffer[4020] = 8'h0c;
 buffer[4021] = 8'h0c;
 buffer[4022] = 8'h0c;
 buffer[4023] = 8'hec;
 buffer[4024] = 8'h6c;
 buffer[4025] = 8'h6c;
 buffer[4026] = 8'h3c;
 buffer[4027] = 8'h1c;
 buffer[4028] = 8'h00;
 buffer[4029] = 8'h00;
 buffer[4030] = 8'h00;
 buffer[4031] = 8'h00;
 buffer[4032] = 8'h00;
 buffer[4033] = 8'hd8;
 buffer[4034] = 8'h6c;
 buffer[4035] = 8'h6c;
 buffer[4036] = 8'h6c;
 buffer[4037] = 8'h6c;
 buffer[4038] = 8'h6c;
 buffer[4039] = 8'h00;
 buffer[4040] = 8'h00;
 buffer[4041] = 8'h00;
 buffer[4042] = 8'h00;
 buffer[4043] = 8'h00;
 buffer[4044] = 8'h00;
 buffer[4045] = 8'h00;
 buffer[4046] = 8'h00;
 buffer[4047] = 8'h00;
 buffer[4048] = 8'h00;
 buffer[4049] = 8'h70;
 buffer[4050] = 8'hd8;
 buffer[4051] = 8'h30;
 buffer[4052] = 8'h60;
 buffer[4053] = 8'hc8;
 buffer[4054] = 8'hf8;
 buffer[4055] = 8'h00;
 buffer[4056] = 8'h00;
 buffer[4057] = 8'h00;
 buffer[4058] = 8'h00;
 buffer[4059] = 8'h00;
 buffer[4060] = 8'h00;
 buffer[4061] = 8'h00;
 buffer[4062] = 8'h00;
 buffer[4063] = 8'h00;
 buffer[4064] = 8'h00;
 buffer[4065] = 8'h00;
 buffer[4066] = 8'h00;
 buffer[4067] = 8'h00;
 buffer[4068] = 8'h7c;
 buffer[4069] = 8'h7c;
 buffer[4070] = 8'h7c;
 buffer[4071] = 8'h7c;
 buffer[4072] = 8'h7c;
 buffer[4073] = 8'h7c;
 buffer[4074] = 8'h7c;
 buffer[4075] = 8'h00;
 buffer[4076] = 8'h00;
 buffer[4077] = 8'h00;
 buffer[4078] = 8'h00;
 buffer[4079] = 8'h00;
 buffer[4080] = 8'h00;
 buffer[4081] = 8'h00;
 buffer[4082] = 8'h00;
 buffer[4083] = 8'h00;
 buffer[4084] = 8'h00;
 buffer[4085] = 8'h00;
 buffer[4086] = 8'h00;
 buffer[4087] = 8'h00;
 buffer[4088] = 8'h00;
 buffer[4089] = 8'h00;
 buffer[4090] = 8'h00;
 buffer[4091] = 8'h00;
 buffer[4092] = 8'h00;
 buffer[4093] = 8'h00;
 buffer[4094] = 8'h00;
 buffer[4095] = 8'h00;
end

endmodule

module M_character_map_mem_charactermap(
input      [11:0]                in_charactermap_addr0,
output reg  [20:0]     out_charactermap_rdata0,
output reg  [20:0]     out_charactermap_rdata1,
input      [0:0]             in_charactermap_wenable1,
input      [20:0]                 in_charactermap_wdata1,
input      [11:0]                in_charactermap_addr1,
input      clock0,
input      clock1
);
reg  [20:0] buffer[2399:0];
always @(posedge clock0) begin
  out_charactermap_rdata0 <= buffer[in_charactermap_addr0];
end
always @(posedge clock1) begin
  if (in_charactermap_wenable1) begin
    buffer[in_charactermap_addr1] <= in_charactermap_wdata1;
  end
end
initial begin
 buffer[0] = 21'b100000000000000000000;
 buffer[1] = 21'b100000000000000000000;
 buffer[2] = 21'b100000000000000000000;
 buffer[3] = 21'b100000000000000000000;
 buffer[4] = 21'b100000000000000000000;
 buffer[5] = 21'b100000000000000000000;
 buffer[6] = 21'b100000000000000000000;
 buffer[7] = 21'b100000000000000000000;
 buffer[8] = 21'b100000000000000000000;
 buffer[9] = 21'b100000000000000000000;
 buffer[10] = 21'b100000000000000000000;
 buffer[11] = 21'b100000000000000000000;
 buffer[12] = 21'b100000000000000000000;
 buffer[13] = 21'b100000000000000000000;
 buffer[14] = 21'b100000000000000000000;
 buffer[15] = 21'b100000000000000000000;
 buffer[16] = 21'b100000000000000000000;
 buffer[17] = 21'b100000000000000000000;
 buffer[18] = 21'b100000000000000000000;
 buffer[19] = 21'b100000000000000000000;
 buffer[20] = 21'b100000000000000000000;
 buffer[21] = 21'b100000000000000000000;
 buffer[22] = 21'b100000000000000000000;
 buffer[23] = 21'b100000000000000000000;
 buffer[24] = 21'b100000000000000000000;
 buffer[25] = 21'b100000000000000000000;
 buffer[26] = 21'b100000000000000000000;
 buffer[27] = 21'b100000000000000000000;
 buffer[28] = 21'b100000000000000000000;
 buffer[29] = 21'b100000000000000000000;
 buffer[30] = 21'b100000000000000000000;
 buffer[31] = 21'b100000000000000000000;
 buffer[32] = 21'b100000000000000000000;
 buffer[33] = 21'b100000000000000000000;
 buffer[34] = 21'b100000000000000000000;
 buffer[35] = 21'b100000000000000000000;
 buffer[36] = 21'b100000000000000000000;
 buffer[37] = 21'b100000000000000000000;
 buffer[38] = 21'b100000000000000000000;
 buffer[39] = 21'b100000000000000000000;
 buffer[40] = 21'b100000000000000000000;
 buffer[41] = 21'b100000000000000000000;
 buffer[42] = 21'b100000000000000000000;
 buffer[43] = 21'b100000000000000000000;
 buffer[44] = 21'b100000000000000000000;
 buffer[45] = 21'b100000000000000000000;
 buffer[46] = 21'b100000000000000000000;
 buffer[47] = 21'b100000000000000000000;
 buffer[48] = 21'b100000000000000000000;
 buffer[49] = 21'b100000000000000000000;
 buffer[50] = 21'b100000000000000000000;
 buffer[51] = 21'b100000000000000000000;
 buffer[52] = 21'b100000000000000000000;
 buffer[53] = 21'b100000000000000000000;
 buffer[54] = 21'b100000000000000000000;
 buffer[55] = 21'b100000000000000000000;
 buffer[56] = 21'b100000000000000000000;
 buffer[57] = 21'b100000000000000000000;
 buffer[58] = 21'b100000000000000000000;
 buffer[59] = 21'b100000000000000000000;
 buffer[60] = 21'b100000000000000000000;
 buffer[61] = 21'b100000000000000000000;
 buffer[62] = 21'b100000000000000000000;
 buffer[63] = 21'b100000000000000000000;
 buffer[64] = 21'b100000000000000000000;
 buffer[65] = 21'b100000000000000000000;
 buffer[66] = 21'b100000000000000000000;
 buffer[67] = 21'b100000000000000000000;
 buffer[68] = 21'b100000000000000000000;
 buffer[69] = 21'b100000000000000000000;
 buffer[70] = 21'b100000000000000000000;
 buffer[71] = 21'b100000000000000000000;
 buffer[72] = 21'b100000000000000000000;
 buffer[73] = 21'b100000000000000000000;
 buffer[74] = 21'b100000000000000000000;
 buffer[75] = 21'b100000000000000000000;
 buffer[76] = 21'b100000000000000000000;
 buffer[77] = 21'b100000000000000000000;
 buffer[78] = 21'b100000000000000000000;
 buffer[79] = 21'b100000000000000000000;
 buffer[80] = 21'b100000000000000000000;
 buffer[81] = 21'b100000000000000000000;
 buffer[82] = 21'b100000000000000000000;
 buffer[83] = 21'b100000000000000000000;
 buffer[84] = 21'b100000000000000000000;
 buffer[85] = 21'b100000000000000000000;
 buffer[86] = 21'b100000000000000000000;
 buffer[87] = 21'b100000000000000000000;
 buffer[88] = 21'b100000000000000000000;
 buffer[89] = 21'b100000000000000000000;
 buffer[90] = 21'b100000000000000000000;
 buffer[91] = 21'b100000000000000000000;
 buffer[92] = 21'b100000000000000000000;
 buffer[93] = 21'b100000000000000000000;
 buffer[94] = 21'b100000000000000000000;
 buffer[95] = 21'b100000000000000000000;
 buffer[96] = 21'b100000000000000000000;
 buffer[97] = 21'b100000000000000000000;
 buffer[98] = 21'b100000000000000000000;
 buffer[99] = 21'b100000000000000000000;
 buffer[100] = 21'b100000000000000000000;
 buffer[101] = 21'b100000000000000000000;
 buffer[102] = 21'b100000000000000000000;
 buffer[103] = 21'b100000000000000000000;
 buffer[104] = 21'b100000000000000000000;
 buffer[105] = 21'b100000000000000000000;
 buffer[106] = 21'b100000000000000000000;
 buffer[107] = 21'b100000000000000000000;
 buffer[108] = 21'b100000000000000000000;
 buffer[109] = 21'b100000000000000000000;
 buffer[110] = 21'b100000000000000000000;
 buffer[111] = 21'b100000000000000000000;
 buffer[112] = 21'b100000000000000000000;
 buffer[113] = 21'b100000000000000000000;
 buffer[114] = 21'b100000000000000000000;
 buffer[115] = 21'b100000000000000000000;
 buffer[116] = 21'b100000000000000000000;
 buffer[117] = 21'b100000000000000000000;
 buffer[118] = 21'b100000000000000000000;
 buffer[119] = 21'b100000000000000000000;
 buffer[120] = 21'b100000000000000000000;
 buffer[121] = 21'b100000000000000000000;
 buffer[122] = 21'b100000000000000000000;
 buffer[123] = 21'b100000000000000000000;
 buffer[124] = 21'b100000000000000000000;
 buffer[125] = 21'b100000000000000000000;
 buffer[126] = 21'b100000000000000000000;
 buffer[127] = 21'b100000000000000000000;
 buffer[128] = 21'b100000000000000000000;
 buffer[129] = 21'b100000000000000000000;
 buffer[130] = 21'b100000000000000000000;
 buffer[131] = 21'b100000000000000000000;
 buffer[132] = 21'b100000000000000000000;
 buffer[133] = 21'b100000000000000000000;
 buffer[134] = 21'b100000000000000000000;
 buffer[135] = 21'b100000000000000000000;
 buffer[136] = 21'b100000000000000000000;
 buffer[137] = 21'b100000000000000000000;
 buffer[138] = 21'b100000000000000000000;
 buffer[139] = 21'b100000000000000000000;
 buffer[140] = 21'b100000000000000000000;
 buffer[141] = 21'b100000000000000000000;
 buffer[142] = 21'b100000000000000000000;
 buffer[143] = 21'b100000000000000000000;
 buffer[144] = 21'b100000000000000000000;
 buffer[145] = 21'b100000000000000000000;
 buffer[146] = 21'b100000000000000000000;
 buffer[147] = 21'b100000000000000000000;
 buffer[148] = 21'b100000000000000000000;
 buffer[149] = 21'b100000000000000000000;
 buffer[150] = 21'b100000000000000000000;
 buffer[151] = 21'b100000000000000000000;
 buffer[152] = 21'b100000000000000000000;
 buffer[153] = 21'b100000000000000000000;
 buffer[154] = 21'b100000000000000000000;
 buffer[155] = 21'b100000000000000000000;
 buffer[156] = 21'b100000000000000000000;
 buffer[157] = 21'b100000000000000000000;
 buffer[158] = 21'b100000000000000000000;
 buffer[159] = 21'b100000000000000000000;
 buffer[160] = 21'b100000000000000000000;
 buffer[161] = 21'b100000000000000000000;
 buffer[162] = 21'b100000000000000000000;
 buffer[163] = 21'b100000000000000000000;
 buffer[164] = 21'b100000000000000000000;
 buffer[165] = 21'b100000000000000000000;
 buffer[166] = 21'b100000000000000000000;
 buffer[167] = 21'b100000000000000000000;
 buffer[168] = 21'b100000000000000000000;
 buffer[169] = 21'b100000000000000000000;
 buffer[170] = 21'b100000000000000000000;
 buffer[171] = 21'b100000000000000000000;
 buffer[172] = 21'b100000000000000000000;
 buffer[173] = 21'b100000000000000000000;
 buffer[174] = 21'b100000000000000000000;
 buffer[175] = 21'b100000000000000000000;
 buffer[176] = 21'b100000000000000000000;
 buffer[177] = 21'b100000000000000000000;
 buffer[178] = 21'b100000000000000000000;
 buffer[179] = 21'b100000000000000000000;
 buffer[180] = 21'b100000000000000000000;
 buffer[181] = 21'b100000000000000000000;
 buffer[182] = 21'b100000000000000000000;
 buffer[183] = 21'b100000000000000000000;
 buffer[184] = 21'b100000000000000000000;
 buffer[185] = 21'b100000000000000000000;
 buffer[186] = 21'b100000000000000000000;
 buffer[187] = 21'b100000000000000000000;
 buffer[188] = 21'b100000000000000000000;
 buffer[189] = 21'b100000000000000000000;
 buffer[190] = 21'b100000000000000000000;
 buffer[191] = 21'b100000000000000000000;
 buffer[192] = 21'b100000000000000000000;
 buffer[193] = 21'b100000000000000000000;
 buffer[194] = 21'b100000000000000000000;
 buffer[195] = 21'b100000000000000000000;
 buffer[196] = 21'b100000000000000000000;
 buffer[197] = 21'b100000000000000000000;
 buffer[198] = 21'b100000000000000000000;
 buffer[199] = 21'b100000000000000000000;
 buffer[200] = 21'b100000000000000000000;
 buffer[201] = 21'b100000000000000000000;
 buffer[202] = 21'b100000000000000000000;
 buffer[203] = 21'b100000000000000000000;
 buffer[204] = 21'b100000000000000000000;
 buffer[205] = 21'b100000000000000000000;
 buffer[206] = 21'b100000000000000000000;
 buffer[207] = 21'b100000000000000000000;
 buffer[208] = 21'b100000000000000000000;
 buffer[209] = 21'b100000000000000000000;
 buffer[210] = 21'b100000000000000000000;
 buffer[211] = 21'b100000000000000000000;
 buffer[212] = 21'b100000000000000000000;
 buffer[213] = 21'b100000000000000000000;
 buffer[214] = 21'b100000000000000000000;
 buffer[215] = 21'b100000000000000000000;
 buffer[216] = 21'b100000000000000000000;
 buffer[217] = 21'b100000000000000000000;
 buffer[218] = 21'b100000000000000000000;
 buffer[219] = 21'b100000000000000000000;
 buffer[220] = 21'b100000000000000000000;
 buffer[221] = 21'b100000000000000000000;
 buffer[222] = 21'b100000000000000000000;
 buffer[223] = 21'b100000000000000000000;
 buffer[224] = 21'b100000000000000000000;
 buffer[225] = 21'b100000000000000000000;
 buffer[226] = 21'b100000000000000000000;
 buffer[227] = 21'b100000000000000000000;
 buffer[228] = 21'b100000000000000000000;
 buffer[229] = 21'b100000000000000000000;
 buffer[230] = 21'b100000000000000000000;
 buffer[231] = 21'b100000000000000000000;
 buffer[232] = 21'b100000000000000000000;
 buffer[233] = 21'b100000000000000000000;
 buffer[234] = 21'b100000000000000000000;
 buffer[235] = 21'b100000000000000000000;
 buffer[236] = 21'b100000000000000000000;
 buffer[237] = 21'b100000000000000000000;
 buffer[238] = 21'b100000000000000000000;
 buffer[239] = 21'b100000000000000000000;
 buffer[240] = 21'b100000000000000000000;
 buffer[241] = 21'b100000000000000000000;
 buffer[242] = 21'b100000000000000000000;
 buffer[243] = 21'b100000000000000000000;
 buffer[244] = 21'b100000000000000000000;
 buffer[245] = 21'b100000000000000000000;
 buffer[246] = 21'b100000000000000000000;
 buffer[247] = 21'b100000000000000000000;
 buffer[248] = 21'b100000000000000000000;
 buffer[249] = 21'b100000000000000000000;
 buffer[250] = 21'b100000000000000000000;
 buffer[251] = 21'b100000000000000000000;
 buffer[252] = 21'b100000000000000000000;
 buffer[253] = 21'b100000000000000000000;
 buffer[254] = 21'b100000000000000000000;
 buffer[255] = 21'b100000000000000000000;
 buffer[256] = 21'b100000000000000000000;
 buffer[257] = 21'b100000000000000000000;
 buffer[258] = 21'b100000000000000000000;
 buffer[259] = 21'b100000000000000000000;
 buffer[260] = 21'b100000000000000000000;
 buffer[261] = 21'b100000000000000000000;
 buffer[262] = 21'b100000000000000000000;
 buffer[263] = 21'b100000000000000000000;
 buffer[264] = 21'b100000000000000000000;
 buffer[265] = 21'b100000000000000000000;
 buffer[266] = 21'b100000000000000000000;
 buffer[267] = 21'b100000000000000000000;
 buffer[268] = 21'b100000000000000000000;
 buffer[269] = 21'b100000000000000000000;
 buffer[270] = 21'b100000000000000000000;
 buffer[271] = 21'b100000000000000000000;
 buffer[272] = 21'b100000000000000000000;
 buffer[273] = 21'b100000000000000000000;
 buffer[274] = 21'b100000000000000000000;
 buffer[275] = 21'b100000000000000000000;
 buffer[276] = 21'b100000000000000000000;
 buffer[277] = 21'b100000000000000000000;
 buffer[278] = 21'b100000000000000000000;
 buffer[279] = 21'b100000000000000000000;
 buffer[280] = 21'b100000000000000000000;
 buffer[281] = 21'b100000000000000000000;
 buffer[282] = 21'b100000000000000000000;
 buffer[283] = 21'b100000000000000000000;
 buffer[284] = 21'b100000000000000000000;
 buffer[285] = 21'b100000000000000000000;
 buffer[286] = 21'b100000000000000000000;
 buffer[287] = 21'b100000000000000000000;
 buffer[288] = 21'b100000000000000000000;
 buffer[289] = 21'b100000000000000000000;
 buffer[290] = 21'b100000000000000000000;
 buffer[291] = 21'b100000000000000000000;
 buffer[292] = 21'b100000000000000000000;
 buffer[293] = 21'b100000000000000000000;
 buffer[294] = 21'b100000000000000000000;
 buffer[295] = 21'b100000000000000000000;
 buffer[296] = 21'b100000000000000000000;
 buffer[297] = 21'b100000000000000000000;
 buffer[298] = 21'b100000000000000000000;
 buffer[299] = 21'b100000000000000000000;
 buffer[300] = 21'b100000000000000000000;
 buffer[301] = 21'b100000000000000000000;
 buffer[302] = 21'b100000000000000000000;
 buffer[303] = 21'b100000000000000000000;
 buffer[304] = 21'b100000000000000000000;
 buffer[305] = 21'b100000000000000000000;
 buffer[306] = 21'b100000000000000000000;
 buffer[307] = 21'b100000000000000000000;
 buffer[308] = 21'b100000000000000000000;
 buffer[309] = 21'b100000000000000000000;
 buffer[310] = 21'b100000000000000000000;
 buffer[311] = 21'b100000000000000000000;
 buffer[312] = 21'b100000000000000000000;
 buffer[313] = 21'b100000000000000000000;
 buffer[314] = 21'b100000000000000000000;
 buffer[315] = 21'b100000000000000000000;
 buffer[316] = 21'b100000000000000000000;
 buffer[317] = 21'b100000000000000000000;
 buffer[318] = 21'b100000000000000000000;
 buffer[319] = 21'b100000000000000000000;
 buffer[320] = 21'b100000000000000000000;
 buffer[321] = 21'b100000000000000000000;
 buffer[322] = 21'b100000000000000000000;
 buffer[323] = 21'b100000000000000000000;
 buffer[324] = 21'b100000000000000000000;
 buffer[325] = 21'b100000000000000000000;
 buffer[326] = 21'b100000000000000000000;
 buffer[327] = 21'b100000000000000000000;
 buffer[328] = 21'b100000000000000000000;
 buffer[329] = 21'b100000000000000000000;
 buffer[330] = 21'b100000000000000000000;
 buffer[331] = 21'b100000000000000000000;
 buffer[332] = 21'b100000000000000000000;
 buffer[333] = 21'b100000000000000000000;
 buffer[334] = 21'b100000000000000000000;
 buffer[335] = 21'b100000000000000000000;
 buffer[336] = 21'b100000000000000000000;
 buffer[337] = 21'b100000000000000000000;
 buffer[338] = 21'b100000000000000000000;
 buffer[339] = 21'b100000000000000000000;
 buffer[340] = 21'b100000000000000000000;
 buffer[341] = 21'b100000000000000000000;
 buffer[342] = 21'b100000000000000000000;
 buffer[343] = 21'b100000000000000000000;
 buffer[344] = 21'b100000000000000000000;
 buffer[345] = 21'b100000000000000000000;
 buffer[346] = 21'b100000000000000000000;
 buffer[347] = 21'b100000000000000000000;
 buffer[348] = 21'b100000000000000000000;
 buffer[349] = 21'b100000000000000000000;
 buffer[350] = 21'b100000000000000000000;
 buffer[351] = 21'b100000000000000000000;
 buffer[352] = 21'b100000000000000000000;
 buffer[353] = 21'b100000000000000000000;
 buffer[354] = 21'b100000000000000000000;
 buffer[355] = 21'b100000000000000000000;
 buffer[356] = 21'b100000000000000000000;
 buffer[357] = 21'b100000000000000000000;
 buffer[358] = 21'b100000000000000000000;
 buffer[359] = 21'b100000000000000000000;
 buffer[360] = 21'b100000000000000000000;
 buffer[361] = 21'b100000000000000000000;
 buffer[362] = 21'b100000000000000000000;
 buffer[363] = 21'b100000000000000000000;
 buffer[364] = 21'b100000000000000000000;
 buffer[365] = 21'b100000000000000000000;
 buffer[366] = 21'b100000000000000000000;
 buffer[367] = 21'b100000000000000000000;
 buffer[368] = 21'b100000000000000000000;
 buffer[369] = 21'b100000000000000000000;
 buffer[370] = 21'b100000000000000000000;
 buffer[371] = 21'b100000000000000000000;
 buffer[372] = 21'b100000000000000000000;
 buffer[373] = 21'b100000000000000000000;
 buffer[374] = 21'b100000000000000000000;
 buffer[375] = 21'b100000000000000000000;
 buffer[376] = 21'b100000000000000000000;
 buffer[377] = 21'b100000000000000000000;
 buffer[378] = 21'b100000000000000000000;
 buffer[379] = 21'b100000000000000000000;
 buffer[380] = 21'b100000000000000000000;
 buffer[381] = 21'b100000000000000000000;
 buffer[382] = 21'b100000000000000000000;
 buffer[383] = 21'b100000000000000000000;
 buffer[384] = 21'b100000000000000000000;
 buffer[385] = 21'b100000000000000000000;
 buffer[386] = 21'b100000000000000000000;
 buffer[387] = 21'b100000000000000000000;
 buffer[388] = 21'b100000000000000000000;
 buffer[389] = 21'b100000000000000000000;
 buffer[390] = 21'b100000000000000000000;
 buffer[391] = 21'b100000000000000000000;
 buffer[392] = 21'b100000000000000000000;
 buffer[393] = 21'b100000000000000000000;
 buffer[394] = 21'b100000000000000000000;
 buffer[395] = 21'b100000000000000000000;
 buffer[396] = 21'b100000000000000000000;
 buffer[397] = 21'b100000000000000000000;
 buffer[398] = 21'b100000000000000000000;
 buffer[399] = 21'b100000000000000000000;
 buffer[400] = 21'b100000000000000000000;
 buffer[401] = 21'b100000000000000000000;
 buffer[402] = 21'b100000000000000000000;
 buffer[403] = 21'b100000000000000000000;
 buffer[404] = 21'b100000000000000000000;
 buffer[405] = 21'b100000000000000000000;
 buffer[406] = 21'b100000000000000000000;
 buffer[407] = 21'b100000000000000000000;
 buffer[408] = 21'b100000000000000000000;
 buffer[409] = 21'b100000000000000000000;
 buffer[410] = 21'b100000000000000000000;
 buffer[411] = 21'b100000000000000000000;
 buffer[412] = 21'b100000000000000000000;
 buffer[413] = 21'b100000000000000000000;
 buffer[414] = 21'b100000000000000000000;
 buffer[415] = 21'b100000000000000000000;
 buffer[416] = 21'b100000000000000000000;
 buffer[417] = 21'b100000000000000000000;
 buffer[418] = 21'b100000000000000000000;
 buffer[419] = 21'b100000000000000000000;
 buffer[420] = 21'b100000000000000000000;
 buffer[421] = 21'b100000000000000000000;
 buffer[422] = 21'b100000000000000000000;
 buffer[423] = 21'b100000000000000000000;
 buffer[424] = 21'b100000000000000000000;
 buffer[425] = 21'b100000000000000000000;
 buffer[426] = 21'b100000000000000000000;
 buffer[427] = 21'b100000000000000000000;
 buffer[428] = 21'b100000000000000000000;
 buffer[429] = 21'b100000000000000000000;
 buffer[430] = 21'b100000000000000000000;
 buffer[431] = 21'b100000000000000000000;
 buffer[432] = 21'b100000000000000000000;
 buffer[433] = 21'b100000000000000000000;
 buffer[434] = 21'b100000000000000000000;
 buffer[435] = 21'b100000000000000000000;
 buffer[436] = 21'b100000000000000000000;
 buffer[437] = 21'b100000000000000000000;
 buffer[438] = 21'b100000000000000000000;
 buffer[439] = 21'b100000000000000000000;
 buffer[440] = 21'b100000000000000000000;
 buffer[441] = 21'b100000000000000000000;
 buffer[442] = 21'b100000000000000000000;
 buffer[443] = 21'b100000000000000000000;
 buffer[444] = 21'b100000000000000000000;
 buffer[445] = 21'b100000000000000000000;
 buffer[446] = 21'b100000000000000000000;
 buffer[447] = 21'b100000000000000000000;
 buffer[448] = 21'b100000000000000000000;
 buffer[449] = 21'b100000000000000000000;
 buffer[450] = 21'b100000000000000000000;
 buffer[451] = 21'b100000000000000000000;
 buffer[452] = 21'b100000000000000000000;
 buffer[453] = 21'b100000000000000000000;
 buffer[454] = 21'b100000000000000000000;
 buffer[455] = 21'b100000000000000000000;
 buffer[456] = 21'b100000000000000000000;
 buffer[457] = 21'b100000000000000000000;
 buffer[458] = 21'b100000000000000000000;
 buffer[459] = 21'b100000000000000000000;
 buffer[460] = 21'b100000000000000000000;
 buffer[461] = 21'b100000000000000000000;
 buffer[462] = 21'b100000000000000000000;
 buffer[463] = 21'b100000000000000000000;
 buffer[464] = 21'b100000000000000000000;
 buffer[465] = 21'b100000000000000000000;
 buffer[466] = 21'b100000000000000000000;
 buffer[467] = 21'b100000000000000000000;
 buffer[468] = 21'b100000000000000000000;
 buffer[469] = 21'b100000000000000000000;
 buffer[470] = 21'b100000000000000000000;
 buffer[471] = 21'b100000000000000000000;
 buffer[472] = 21'b100000000000000000000;
 buffer[473] = 21'b100000000000000000000;
 buffer[474] = 21'b100000000000000000000;
 buffer[475] = 21'b100000000000000000000;
 buffer[476] = 21'b100000000000000000000;
 buffer[477] = 21'b100000000000000000000;
 buffer[478] = 21'b100000000000000000000;
 buffer[479] = 21'b100000000000000000000;
 buffer[480] = 21'b100000000000000000000;
 buffer[481] = 21'b100000000000000000000;
 buffer[482] = 21'b100000000000000000000;
 buffer[483] = 21'b100000000000000000000;
 buffer[484] = 21'b100000000000000000000;
 buffer[485] = 21'b100000000000000000000;
 buffer[486] = 21'b100000000000000000000;
 buffer[487] = 21'b100000000000000000000;
 buffer[488] = 21'b100000000000000000000;
 buffer[489] = 21'b100000000000000000000;
 buffer[490] = 21'b100000000000000000000;
 buffer[491] = 21'b100000000000000000000;
 buffer[492] = 21'b100000000000000000000;
 buffer[493] = 21'b100000000000000000000;
 buffer[494] = 21'b100000000000000000000;
 buffer[495] = 21'b100000000000000000000;
 buffer[496] = 21'b100000000000000000000;
 buffer[497] = 21'b100000000000000000000;
 buffer[498] = 21'b100000000000000000000;
 buffer[499] = 21'b100000000000000000000;
 buffer[500] = 21'b100000000000000000000;
 buffer[501] = 21'b100000000000000000000;
 buffer[502] = 21'b100000000000000000000;
 buffer[503] = 21'b100000000000000000000;
 buffer[504] = 21'b100000000000000000000;
 buffer[505] = 21'b100000000000000000000;
 buffer[506] = 21'b100000000000000000000;
 buffer[507] = 21'b100000000000000000000;
 buffer[508] = 21'b100000000000000000000;
 buffer[509] = 21'b100000000000000000000;
 buffer[510] = 21'b100000000000000000000;
 buffer[511] = 21'b100000000000000000000;
 buffer[512] = 21'b100000000000000000000;
 buffer[513] = 21'b100000000000000000000;
 buffer[514] = 21'b100000000000000000000;
 buffer[515] = 21'b100000000000000000000;
 buffer[516] = 21'b100000000000000000000;
 buffer[517] = 21'b100000000000000000000;
 buffer[518] = 21'b100000000000000000000;
 buffer[519] = 21'b100000000000000000000;
 buffer[520] = 21'b100000000000000000000;
 buffer[521] = 21'b100000000000000000000;
 buffer[522] = 21'b100000000000000000000;
 buffer[523] = 21'b100000000000000000000;
 buffer[524] = 21'b100000000000000000000;
 buffer[525] = 21'b100000000000000000000;
 buffer[526] = 21'b100000000000000000000;
 buffer[527] = 21'b100000000000000000000;
 buffer[528] = 21'b100000000000000000000;
 buffer[529] = 21'b100000000000000000000;
 buffer[530] = 21'b100000000000000000000;
 buffer[531] = 21'b100000000000000000000;
 buffer[532] = 21'b100000000000000000000;
 buffer[533] = 21'b100000000000000000000;
 buffer[534] = 21'b100000000000000000000;
 buffer[535] = 21'b100000000000000000000;
 buffer[536] = 21'b100000000000000000000;
 buffer[537] = 21'b100000000000000000000;
 buffer[538] = 21'b100000000000000000000;
 buffer[539] = 21'b100000000000000000000;
 buffer[540] = 21'b100000000000000000000;
 buffer[541] = 21'b100000000000000000000;
 buffer[542] = 21'b100000000000000000000;
 buffer[543] = 21'b100000000000000000000;
 buffer[544] = 21'b100000000000000000000;
 buffer[545] = 21'b100000000000000000000;
 buffer[546] = 21'b100000000000000000000;
 buffer[547] = 21'b100000000000000000000;
 buffer[548] = 21'b100000000000000000000;
 buffer[549] = 21'b100000000000000000000;
 buffer[550] = 21'b100000000000000000000;
 buffer[551] = 21'b100000000000000000000;
 buffer[552] = 21'b100000000000000000000;
 buffer[553] = 21'b100000000000000000000;
 buffer[554] = 21'b100000000000000000000;
 buffer[555] = 21'b100000000000000000000;
 buffer[556] = 21'b100000000000000000000;
 buffer[557] = 21'b100000000000000000000;
 buffer[558] = 21'b100000000000000000000;
 buffer[559] = 21'b100000000000000000000;
 buffer[560] = 21'b100000000000000000000;
 buffer[561] = 21'b100000000000000000000;
 buffer[562] = 21'b100000000000000000000;
 buffer[563] = 21'b100000000000000000000;
 buffer[564] = 21'b100000000000000000000;
 buffer[565] = 21'b100000000000000000000;
 buffer[566] = 21'b100000000000000000000;
 buffer[567] = 21'b100000000000000000000;
 buffer[568] = 21'b100000000000000000000;
 buffer[569] = 21'b100000000000000000000;
 buffer[570] = 21'b100000000000000000000;
 buffer[571] = 21'b100000000000000000000;
 buffer[572] = 21'b100000000000000000000;
 buffer[573] = 21'b100000000000000000000;
 buffer[574] = 21'b100000000000000000000;
 buffer[575] = 21'b100000000000000000000;
 buffer[576] = 21'b100000000000000000000;
 buffer[577] = 21'b100000000000000000000;
 buffer[578] = 21'b100000000000000000000;
 buffer[579] = 21'b100000000000000000000;
 buffer[580] = 21'b100000000000000000000;
 buffer[581] = 21'b100000000000000000000;
 buffer[582] = 21'b100000000000000000000;
 buffer[583] = 21'b100000000000000000000;
 buffer[584] = 21'b100000000000000000000;
 buffer[585] = 21'b100000000000000000000;
 buffer[586] = 21'b100000000000000000000;
 buffer[587] = 21'b100000000000000000000;
 buffer[588] = 21'b100000000000000000000;
 buffer[589] = 21'b100000000000000000000;
 buffer[590] = 21'b100000000000000000000;
 buffer[591] = 21'b100000000000000000000;
 buffer[592] = 21'b100000000000000000000;
 buffer[593] = 21'b100000000000000000000;
 buffer[594] = 21'b100000000000000000000;
 buffer[595] = 21'b100000000000000000000;
 buffer[596] = 21'b100000000000000000000;
 buffer[597] = 21'b100000000000000000000;
 buffer[598] = 21'b100000000000000000000;
 buffer[599] = 21'b100000000000000000000;
 buffer[600] = 21'b100000000000000000000;
 buffer[601] = 21'b100000000000000000000;
 buffer[602] = 21'b100000000000000000000;
 buffer[603] = 21'b100000000000000000000;
 buffer[604] = 21'b100000000000000000000;
 buffer[605] = 21'b100000000000000000000;
 buffer[606] = 21'b100000000000000000000;
 buffer[607] = 21'b100000000000000000000;
 buffer[608] = 21'b100000000000000000000;
 buffer[609] = 21'b100000000000000000000;
 buffer[610] = 21'b100000000000000000000;
 buffer[611] = 21'b100000000000000000000;
 buffer[612] = 21'b100000000000000000000;
 buffer[613] = 21'b100000000000000000000;
 buffer[614] = 21'b100000000000000000000;
 buffer[615] = 21'b100000000000000000000;
 buffer[616] = 21'b100000000000000000000;
 buffer[617] = 21'b100000000000000000000;
 buffer[618] = 21'b100000000000000000000;
 buffer[619] = 21'b100000000000000000000;
 buffer[620] = 21'b100000000000000000000;
 buffer[621] = 21'b100000000000000000000;
 buffer[622] = 21'b100000000000000000000;
 buffer[623] = 21'b100000000000000000000;
 buffer[624] = 21'b100000000000000000000;
 buffer[625] = 21'b100000000000000000000;
 buffer[626] = 21'b100000000000000000000;
 buffer[627] = 21'b100000000000000000000;
 buffer[628] = 21'b100000000000000000000;
 buffer[629] = 21'b100000000000000000000;
 buffer[630] = 21'b100000000000000000000;
 buffer[631] = 21'b100000000000000000000;
 buffer[632] = 21'b100000000000000000000;
 buffer[633] = 21'b100000000000000000000;
 buffer[634] = 21'b100000000000000000000;
 buffer[635] = 21'b100000000000000000000;
 buffer[636] = 21'b100000000000000000000;
 buffer[637] = 21'b100000000000000000000;
 buffer[638] = 21'b100000000000000000000;
 buffer[639] = 21'b100000000000000000000;
 buffer[640] = 21'b100000000000000000000;
 buffer[641] = 21'b100000000000000000000;
 buffer[642] = 21'b100000000000000000000;
 buffer[643] = 21'b100000000000000000000;
 buffer[644] = 21'b100000000000000000000;
 buffer[645] = 21'b100000000000000000000;
 buffer[646] = 21'b100000000000000000000;
 buffer[647] = 21'b100000000000000000000;
 buffer[648] = 21'b100000000000000000000;
 buffer[649] = 21'b100000000000000000000;
 buffer[650] = 21'b100000000000000000000;
 buffer[651] = 21'b100000000000000000000;
 buffer[652] = 21'b100000000000000000000;
 buffer[653] = 21'b100000000000000000000;
 buffer[654] = 21'b100000000000000000000;
 buffer[655] = 21'b100000000000000000000;
 buffer[656] = 21'b100000000000000000000;
 buffer[657] = 21'b100000000000000000000;
 buffer[658] = 21'b100000000000000000000;
 buffer[659] = 21'b100000000000000000000;
 buffer[660] = 21'b100000000000000000000;
 buffer[661] = 21'b100000000000000000000;
 buffer[662] = 21'b100000000000000000000;
 buffer[663] = 21'b100000000000000000000;
 buffer[664] = 21'b100000000000000000000;
 buffer[665] = 21'b100000000000000000000;
 buffer[666] = 21'b100000000000000000000;
 buffer[667] = 21'b100000000000000000000;
 buffer[668] = 21'b100000000000000000000;
 buffer[669] = 21'b100000000000000000000;
 buffer[670] = 21'b100000000000000000000;
 buffer[671] = 21'b100000000000000000000;
 buffer[672] = 21'b100000000000000000000;
 buffer[673] = 21'b100000000000000000000;
 buffer[674] = 21'b100000000000000000000;
 buffer[675] = 21'b100000000000000000000;
 buffer[676] = 21'b100000000000000000000;
 buffer[677] = 21'b100000000000000000000;
 buffer[678] = 21'b100000000000000000000;
 buffer[679] = 21'b100000000000000000000;
 buffer[680] = 21'b100000000000000000000;
 buffer[681] = 21'b100000000000000000000;
 buffer[682] = 21'b100000000000000000000;
 buffer[683] = 21'b100000000000000000000;
 buffer[684] = 21'b100000000000000000000;
 buffer[685] = 21'b100000000000000000000;
 buffer[686] = 21'b100000000000000000000;
 buffer[687] = 21'b100000000000000000000;
 buffer[688] = 21'b100000000000000000000;
 buffer[689] = 21'b100000000000000000000;
 buffer[690] = 21'b100000000000000000000;
 buffer[691] = 21'b100000000000000000000;
 buffer[692] = 21'b100000000000000000000;
 buffer[693] = 21'b100000000000000000000;
 buffer[694] = 21'b100000000000000000000;
 buffer[695] = 21'b100000000000000000000;
 buffer[696] = 21'b100000000000000000000;
 buffer[697] = 21'b100000000000000000000;
 buffer[698] = 21'b100000000000000000000;
 buffer[699] = 21'b100000000000000000000;
 buffer[700] = 21'b100000000000000000000;
 buffer[701] = 21'b100000000000000000000;
 buffer[702] = 21'b100000000000000000000;
 buffer[703] = 21'b100000000000000000000;
 buffer[704] = 21'b100000000000000000000;
 buffer[705] = 21'b100000000000000000000;
 buffer[706] = 21'b100000000000000000000;
 buffer[707] = 21'b100000000000000000000;
 buffer[708] = 21'b100000000000000000000;
 buffer[709] = 21'b100000000000000000000;
 buffer[710] = 21'b100000000000000000000;
 buffer[711] = 21'b100000000000000000000;
 buffer[712] = 21'b100000000000000000000;
 buffer[713] = 21'b100000000000000000000;
 buffer[714] = 21'b100000000000000000000;
 buffer[715] = 21'b100000000000000000000;
 buffer[716] = 21'b100000000000000000000;
 buffer[717] = 21'b100000000000000000000;
 buffer[718] = 21'b100000000000000000000;
 buffer[719] = 21'b100000000000000000000;
 buffer[720] = 21'b100000000000000000000;
 buffer[721] = 21'b100000000000000000000;
 buffer[722] = 21'b100000000000000000000;
 buffer[723] = 21'b100000000000000000000;
 buffer[724] = 21'b100000000000000000000;
 buffer[725] = 21'b100000000000000000000;
 buffer[726] = 21'b100000000000000000000;
 buffer[727] = 21'b100000000000000000000;
 buffer[728] = 21'b100000000000000000000;
 buffer[729] = 21'b100000000000000000000;
 buffer[730] = 21'b100000000000000000000;
 buffer[731] = 21'b100000000000000000000;
 buffer[732] = 21'b100000000000000000000;
 buffer[733] = 21'b100000000000000000000;
 buffer[734] = 21'b100000000000000000000;
 buffer[735] = 21'b100000000000000000000;
 buffer[736] = 21'b100000000000000000000;
 buffer[737] = 21'b100000000000000000000;
 buffer[738] = 21'b100000000000000000000;
 buffer[739] = 21'b100000000000000000000;
 buffer[740] = 21'b100000000000000000000;
 buffer[741] = 21'b100000000000000000000;
 buffer[742] = 21'b100000000000000000000;
 buffer[743] = 21'b100000000000000000000;
 buffer[744] = 21'b100000000000000000000;
 buffer[745] = 21'b100000000000000000000;
 buffer[746] = 21'b100000000000000000000;
 buffer[747] = 21'b100000000000000000000;
 buffer[748] = 21'b100000000000000000000;
 buffer[749] = 21'b100000000000000000000;
 buffer[750] = 21'b100000000000000000000;
 buffer[751] = 21'b100000000000000000000;
 buffer[752] = 21'b100000000000000000000;
 buffer[753] = 21'b100000000000000000000;
 buffer[754] = 21'b100000000000000000000;
 buffer[755] = 21'b100000000000000000000;
 buffer[756] = 21'b100000000000000000000;
 buffer[757] = 21'b100000000000000000000;
 buffer[758] = 21'b100000000000000000000;
 buffer[759] = 21'b100000000000000000000;
 buffer[760] = 21'b100000000000000000000;
 buffer[761] = 21'b100000000000000000000;
 buffer[762] = 21'b100000000000000000000;
 buffer[763] = 21'b100000000000000000000;
 buffer[764] = 21'b100000000000000000000;
 buffer[765] = 21'b100000000000000000000;
 buffer[766] = 21'b100000000000000000000;
 buffer[767] = 21'b100000000000000000000;
 buffer[768] = 21'b100000000000000000000;
 buffer[769] = 21'b100000000000000000000;
 buffer[770] = 21'b100000000000000000000;
 buffer[771] = 21'b100000000000000000000;
 buffer[772] = 21'b100000000000000000000;
 buffer[773] = 21'b100000000000000000000;
 buffer[774] = 21'b100000000000000000000;
 buffer[775] = 21'b100000000000000000000;
 buffer[776] = 21'b100000000000000000000;
 buffer[777] = 21'b100000000000000000000;
 buffer[778] = 21'b100000000000000000000;
 buffer[779] = 21'b100000000000000000000;
 buffer[780] = 21'b100000000000000000000;
 buffer[781] = 21'b100000000000000000000;
 buffer[782] = 21'b100000000000000000000;
 buffer[783] = 21'b100000000000000000000;
 buffer[784] = 21'b100000000000000000000;
 buffer[785] = 21'b100000000000000000000;
 buffer[786] = 21'b100000000000000000000;
 buffer[787] = 21'b100000000000000000000;
 buffer[788] = 21'b100000000000000000000;
 buffer[789] = 21'b100000000000000000000;
 buffer[790] = 21'b100000000000000000000;
 buffer[791] = 21'b100000000000000000000;
 buffer[792] = 21'b100000000000000000000;
 buffer[793] = 21'b100000000000000000000;
 buffer[794] = 21'b100000000000000000000;
 buffer[795] = 21'b100000000000000000000;
 buffer[796] = 21'b100000000000000000000;
 buffer[797] = 21'b100000000000000000000;
 buffer[798] = 21'b100000000000000000000;
 buffer[799] = 21'b100000000000000000000;
 buffer[800] = 21'b100000000000000000000;
 buffer[801] = 21'b100000000000000000000;
 buffer[802] = 21'b100000000000000000000;
 buffer[803] = 21'b100000000000000000000;
 buffer[804] = 21'b100000000000000000000;
 buffer[805] = 21'b100000000000000000000;
 buffer[806] = 21'b100000000000000000000;
 buffer[807] = 21'b100000000000000000000;
 buffer[808] = 21'b100000000000000000000;
 buffer[809] = 21'b100000000000000000000;
 buffer[810] = 21'b100000000000000000000;
 buffer[811] = 21'b100000000000000000000;
 buffer[812] = 21'b100000000000000000000;
 buffer[813] = 21'b100000000000000000000;
 buffer[814] = 21'b100000000000000000000;
 buffer[815] = 21'b100000000000000000000;
 buffer[816] = 21'b100000000000000000000;
 buffer[817] = 21'b100000000000000000000;
 buffer[818] = 21'b100000000000000000000;
 buffer[819] = 21'b100000000000000000000;
 buffer[820] = 21'b100000000000000000000;
 buffer[821] = 21'b100000000000000000000;
 buffer[822] = 21'b100000000000000000000;
 buffer[823] = 21'b100000000000000000000;
 buffer[824] = 21'b100000000000000000000;
 buffer[825] = 21'b100000000000000000000;
 buffer[826] = 21'b100000000000000000000;
 buffer[827] = 21'b100000000000000000000;
 buffer[828] = 21'b100000000000000000000;
 buffer[829] = 21'b100000000000000000000;
 buffer[830] = 21'b100000000000000000000;
 buffer[831] = 21'b100000000000000000000;
 buffer[832] = 21'b100000000000000000000;
 buffer[833] = 21'b100000000000000000000;
 buffer[834] = 21'b100000000000000000000;
 buffer[835] = 21'b100000000000000000000;
 buffer[836] = 21'b100000000000000000000;
 buffer[837] = 21'b100000000000000000000;
 buffer[838] = 21'b100000000000000000000;
 buffer[839] = 21'b100000000000000000000;
 buffer[840] = 21'b100000000000000000000;
 buffer[841] = 21'b100000000000000000000;
 buffer[842] = 21'b100000000000000000000;
 buffer[843] = 21'b100000000000000000000;
 buffer[844] = 21'b100000000000000000000;
 buffer[845] = 21'b100000000000000000000;
 buffer[846] = 21'b100000000000000000000;
 buffer[847] = 21'b100000000000000000000;
 buffer[848] = 21'b100000000000000000000;
 buffer[849] = 21'b100000000000000000000;
 buffer[850] = 21'b100000000000000000000;
 buffer[851] = 21'b100000000000000000000;
 buffer[852] = 21'b100000000000000000000;
 buffer[853] = 21'b100000000000000000000;
 buffer[854] = 21'b100000000000000000000;
 buffer[855] = 21'b100000000000000000000;
 buffer[856] = 21'b100000000000000000000;
 buffer[857] = 21'b100000000000000000000;
 buffer[858] = 21'b100000000000000000000;
 buffer[859] = 21'b100000000000000000000;
 buffer[860] = 21'b100000000000000000000;
 buffer[861] = 21'b100000000000000000000;
 buffer[862] = 21'b100000000000000000000;
 buffer[863] = 21'b100000000000000000000;
 buffer[864] = 21'b100000000000000000000;
 buffer[865] = 21'b100000000000000000000;
 buffer[866] = 21'b100000000000000000000;
 buffer[867] = 21'b100000000000000000000;
 buffer[868] = 21'b100000000000000000000;
 buffer[869] = 21'b100000000000000000000;
 buffer[870] = 21'b100000000000000000000;
 buffer[871] = 21'b100000000000000000000;
 buffer[872] = 21'b100000000000000000000;
 buffer[873] = 21'b100000000000000000000;
 buffer[874] = 21'b100000000000000000000;
 buffer[875] = 21'b100000000000000000000;
 buffer[876] = 21'b100000000000000000000;
 buffer[877] = 21'b100000000000000000000;
 buffer[878] = 21'b100000000000000000000;
 buffer[879] = 21'b100000000000000000000;
 buffer[880] = 21'b100000000000000000000;
 buffer[881] = 21'b100000000000000000000;
 buffer[882] = 21'b100000000000000000000;
 buffer[883] = 21'b100000000000000000000;
 buffer[884] = 21'b100000000000000000000;
 buffer[885] = 21'b100000000000000000000;
 buffer[886] = 21'b100000000000000000000;
 buffer[887] = 21'b100000000000000000000;
 buffer[888] = 21'b100000000000000000000;
 buffer[889] = 21'b100000000000000000000;
 buffer[890] = 21'b100000000000000000000;
 buffer[891] = 21'b100000000000000000000;
 buffer[892] = 21'b100000000000000000000;
 buffer[893] = 21'b100000000000000000000;
 buffer[894] = 21'b100000000000000000000;
 buffer[895] = 21'b100000000000000000000;
 buffer[896] = 21'b100000000000000000000;
 buffer[897] = 21'b100000000000000000000;
 buffer[898] = 21'b100000000000000000000;
 buffer[899] = 21'b100000000000000000000;
 buffer[900] = 21'b100000000000000000000;
 buffer[901] = 21'b100000000000000000000;
 buffer[902] = 21'b100000000000000000000;
 buffer[903] = 21'b100000000000000000000;
 buffer[904] = 21'b100000000000000000000;
 buffer[905] = 21'b100000000000000000000;
 buffer[906] = 21'b100000000000000000000;
 buffer[907] = 21'b100000000000000000000;
 buffer[908] = 21'b100000000000000000000;
 buffer[909] = 21'b100000000000000000000;
 buffer[910] = 21'b100000000000000000000;
 buffer[911] = 21'b100000000000000000000;
 buffer[912] = 21'b100000000000000000000;
 buffer[913] = 21'b100000000000000000000;
 buffer[914] = 21'b100000000000000000000;
 buffer[915] = 21'b100000000000000000000;
 buffer[916] = 21'b100000000000000000000;
 buffer[917] = 21'b100000000000000000000;
 buffer[918] = 21'b100000000000000000000;
 buffer[919] = 21'b100000000000000000000;
 buffer[920] = 21'b100000000000000000000;
 buffer[921] = 21'b100000000000000000000;
 buffer[922] = 21'b100000000000000000000;
 buffer[923] = 21'b100000000000000000000;
 buffer[924] = 21'b100000000000000000000;
 buffer[925] = 21'b100000000000000000000;
 buffer[926] = 21'b100000000000000000000;
 buffer[927] = 21'b100000000000000000000;
 buffer[928] = 21'b100000000000000000000;
 buffer[929] = 21'b100000000000000000000;
 buffer[930] = 21'b100000000000000000000;
 buffer[931] = 21'b100000000000000000000;
 buffer[932] = 21'b100000000000000000000;
 buffer[933] = 21'b100000000000000000000;
 buffer[934] = 21'b100000000000000000000;
 buffer[935] = 21'b100000000000000000000;
 buffer[936] = 21'b100000000000000000000;
 buffer[937] = 21'b100000000000000000000;
 buffer[938] = 21'b100000000000000000000;
 buffer[939] = 21'b100000000000000000000;
 buffer[940] = 21'b100000000000000000000;
 buffer[941] = 21'b100000000000000000000;
 buffer[942] = 21'b100000000000000000000;
 buffer[943] = 21'b100000000000000000000;
 buffer[944] = 21'b100000000000000000000;
 buffer[945] = 21'b100000000000000000000;
 buffer[946] = 21'b100000000000000000000;
 buffer[947] = 21'b100000000000000000000;
 buffer[948] = 21'b100000000000000000000;
 buffer[949] = 21'b100000000000000000000;
 buffer[950] = 21'b100000000000000000000;
 buffer[951] = 21'b100000000000000000000;
 buffer[952] = 21'b100000000000000000000;
 buffer[953] = 21'b100000000000000000000;
 buffer[954] = 21'b100000000000000000000;
 buffer[955] = 21'b100000000000000000000;
 buffer[956] = 21'b100000000000000000000;
 buffer[957] = 21'b100000000000000000000;
 buffer[958] = 21'b100000000000000000000;
 buffer[959] = 21'b100000000000000000000;
 buffer[960] = 21'b100000000000000000000;
 buffer[961] = 21'b100000000000000000000;
 buffer[962] = 21'b100000000000000000000;
 buffer[963] = 21'b100000000000000000000;
 buffer[964] = 21'b100000000000000000000;
 buffer[965] = 21'b100000000000000000000;
 buffer[966] = 21'b100000000000000000000;
 buffer[967] = 21'b100000000000000000000;
 buffer[968] = 21'b100000000000000000000;
 buffer[969] = 21'b100000000000000000000;
 buffer[970] = 21'b100000000000000000000;
 buffer[971] = 21'b100000000000000000000;
 buffer[972] = 21'b100000000000000000000;
 buffer[973] = 21'b100000000000000000000;
 buffer[974] = 21'b100000000000000000000;
 buffer[975] = 21'b100000000000000000000;
 buffer[976] = 21'b100000000000000000000;
 buffer[977] = 21'b100000000000000000000;
 buffer[978] = 21'b100000000000000000000;
 buffer[979] = 21'b100000000000000000000;
 buffer[980] = 21'b100000000000000000000;
 buffer[981] = 21'b100000000000000000000;
 buffer[982] = 21'b100000000000000000000;
 buffer[983] = 21'b100000000000000000000;
 buffer[984] = 21'b100000000000000000000;
 buffer[985] = 21'b100000000000000000000;
 buffer[986] = 21'b100000000000000000000;
 buffer[987] = 21'b100000000000000000000;
 buffer[988] = 21'b100000000000000000000;
 buffer[989] = 21'b100000000000000000000;
 buffer[990] = 21'b100000000000000000000;
 buffer[991] = 21'b100000000000000000000;
 buffer[992] = 21'b100000000000000000000;
 buffer[993] = 21'b100000000000000000000;
 buffer[994] = 21'b100000000000000000000;
 buffer[995] = 21'b100000000000000000000;
 buffer[996] = 21'b100000000000000000000;
 buffer[997] = 21'b100000000000000000000;
 buffer[998] = 21'b100000000000000000000;
 buffer[999] = 21'b100000000000000000000;
 buffer[1000] = 21'b100000000000000000000;
 buffer[1001] = 21'b100000000000000000000;
 buffer[1002] = 21'b100000000000000000000;
 buffer[1003] = 21'b100000000000000000000;
 buffer[1004] = 21'b100000000000000000000;
 buffer[1005] = 21'b100000000000000000000;
 buffer[1006] = 21'b100000000000000000000;
 buffer[1007] = 21'b100000000000000000000;
 buffer[1008] = 21'b100000000000000000000;
 buffer[1009] = 21'b100000000000000000000;
 buffer[1010] = 21'b100000000000000000000;
 buffer[1011] = 21'b100000000000000000000;
 buffer[1012] = 21'b100000000000000000000;
 buffer[1013] = 21'b100000000000000000000;
 buffer[1014] = 21'b100000000000000000000;
 buffer[1015] = 21'b100000000000000000000;
 buffer[1016] = 21'b100000000000000000000;
 buffer[1017] = 21'b100000000000000000000;
 buffer[1018] = 21'b100000000000000000000;
 buffer[1019] = 21'b100000000000000000000;
 buffer[1020] = 21'b100000000000000000000;
 buffer[1021] = 21'b100000000000000000000;
 buffer[1022] = 21'b100000000000000000000;
 buffer[1023] = 21'b100000000000000000000;
 buffer[1024] = 21'b100000000000000000000;
 buffer[1025] = 21'b100000000000000000000;
 buffer[1026] = 21'b100000000000000000000;
 buffer[1027] = 21'b100000000000000000000;
 buffer[1028] = 21'b100000000000000000000;
 buffer[1029] = 21'b100000000000000000000;
 buffer[1030] = 21'b100000000000000000000;
 buffer[1031] = 21'b100000000000000000000;
 buffer[1032] = 21'b100000000000000000000;
 buffer[1033] = 21'b100000000000000000000;
 buffer[1034] = 21'b100000000000000000000;
 buffer[1035] = 21'b100000000000000000000;
 buffer[1036] = 21'b100000000000000000000;
 buffer[1037] = 21'b100000000000000000000;
 buffer[1038] = 21'b100000000000000000000;
 buffer[1039] = 21'b100000000000000000000;
 buffer[1040] = 21'b100000000000000000000;
 buffer[1041] = 21'b100000000000000000000;
 buffer[1042] = 21'b100000000000000000000;
 buffer[1043] = 21'b100000000000000000000;
 buffer[1044] = 21'b100000000000000000000;
 buffer[1045] = 21'b100000000000000000000;
 buffer[1046] = 21'b100000000000000000000;
 buffer[1047] = 21'b100000000000000000000;
 buffer[1048] = 21'b100000000000000000000;
 buffer[1049] = 21'b100000000000000000000;
 buffer[1050] = 21'b100000000000000000000;
 buffer[1051] = 21'b100000000000000000000;
 buffer[1052] = 21'b100000000000000000000;
 buffer[1053] = 21'b100000000000000000000;
 buffer[1054] = 21'b100000000000000000000;
 buffer[1055] = 21'b100000000000000000000;
 buffer[1056] = 21'b100000000000000000000;
 buffer[1057] = 21'b100000000000000000000;
 buffer[1058] = 21'b100000000000000000000;
 buffer[1059] = 21'b100000000000000000000;
 buffer[1060] = 21'b100000000000000000000;
 buffer[1061] = 21'b100000000000000000000;
 buffer[1062] = 21'b100000000000000000000;
 buffer[1063] = 21'b100000000000000000000;
 buffer[1064] = 21'b100000000000000000000;
 buffer[1065] = 21'b100000000000000000000;
 buffer[1066] = 21'b100000000000000000000;
 buffer[1067] = 21'b100000000000000000000;
 buffer[1068] = 21'b100000000000000000000;
 buffer[1069] = 21'b100000000000000000000;
 buffer[1070] = 21'b100000000000000000000;
 buffer[1071] = 21'b100000000000000000000;
 buffer[1072] = 21'b100000000000000000000;
 buffer[1073] = 21'b100000000000000000000;
 buffer[1074] = 21'b100000000000000000000;
 buffer[1075] = 21'b100000000000000000000;
 buffer[1076] = 21'b100000000000000000000;
 buffer[1077] = 21'b100000000000000000000;
 buffer[1078] = 21'b100000000000000000000;
 buffer[1079] = 21'b100000000000000000000;
 buffer[1080] = 21'b100000000000000000000;
 buffer[1081] = 21'b100000000000000000000;
 buffer[1082] = 21'b100000000000000000000;
 buffer[1083] = 21'b100000000000000000000;
 buffer[1084] = 21'b100000000000000000000;
 buffer[1085] = 21'b100000000000000000000;
 buffer[1086] = 21'b100000000000000000000;
 buffer[1087] = 21'b100000000000000000000;
 buffer[1088] = 21'b100000000000000000000;
 buffer[1089] = 21'b100000000000000000000;
 buffer[1090] = 21'b100000000000000000000;
 buffer[1091] = 21'b100000000000000000000;
 buffer[1092] = 21'b100000000000000000000;
 buffer[1093] = 21'b100000000000000000000;
 buffer[1094] = 21'b100000000000000000000;
 buffer[1095] = 21'b100000000000000000000;
 buffer[1096] = 21'b100000000000000000000;
 buffer[1097] = 21'b100000000000000000000;
 buffer[1098] = 21'b100000000000000000000;
 buffer[1099] = 21'b100000000000000000000;
 buffer[1100] = 21'b100000000000000000000;
 buffer[1101] = 21'b100000000000000000000;
 buffer[1102] = 21'b100000000000000000000;
 buffer[1103] = 21'b100000000000000000000;
 buffer[1104] = 21'b100000000000000000000;
 buffer[1105] = 21'b100000000000000000000;
 buffer[1106] = 21'b100000000000000000000;
 buffer[1107] = 21'b100000000000000000000;
 buffer[1108] = 21'b100000000000000000000;
 buffer[1109] = 21'b100000000000000000000;
 buffer[1110] = 21'b100000000000000000000;
 buffer[1111] = 21'b100000000000000000000;
 buffer[1112] = 21'b100000000000000000000;
 buffer[1113] = 21'b100000000000000000000;
 buffer[1114] = 21'b100000000000000000000;
 buffer[1115] = 21'b100000000000000000000;
 buffer[1116] = 21'b100000000000000000000;
 buffer[1117] = 21'b100000000000000000000;
 buffer[1118] = 21'b100000000000000000000;
 buffer[1119] = 21'b100000000000000000000;
 buffer[1120] = 21'b100000000000000000000;
 buffer[1121] = 21'b100000000000000000000;
 buffer[1122] = 21'b100000000000000000000;
 buffer[1123] = 21'b100000000000000000000;
 buffer[1124] = 21'b100000000000000000000;
 buffer[1125] = 21'b100000000000000000000;
 buffer[1126] = 21'b100000000000000000000;
 buffer[1127] = 21'b100000000000000000000;
 buffer[1128] = 21'b100000000000000000000;
 buffer[1129] = 21'b100000000000000000000;
 buffer[1130] = 21'b100000000000000000000;
 buffer[1131] = 21'b100000000000000000000;
 buffer[1132] = 21'b100000000000000000000;
 buffer[1133] = 21'b100000000000000000000;
 buffer[1134] = 21'b100000000000000000000;
 buffer[1135] = 21'b100000000000000000000;
 buffer[1136] = 21'b100000000000000000000;
 buffer[1137] = 21'b100000000000000000000;
 buffer[1138] = 21'b100000000000000000000;
 buffer[1139] = 21'b100000000000000000000;
 buffer[1140] = 21'b100000000000000000000;
 buffer[1141] = 21'b100000000000000000000;
 buffer[1142] = 21'b100000000000000000000;
 buffer[1143] = 21'b100000000000000000000;
 buffer[1144] = 21'b100000000000000000000;
 buffer[1145] = 21'b100000000000000000000;
 buffer[1146] = 21'b100000000000000000000;
 buffer[1147] = 21'b100000000000000000000;
 buffer[1148] = 21'b100000000000000000000;
 buffer[1149] = 21'b100000000000000000000;
 buffer[1150] = 21'b100000000000000000000;
 buffer[1151] = 21'b100000000000000000000;
 buffer[1152] = 21'b100000000000000000000;
 buffer[1153] = 21'b100000000000000000000;
 buffer[1154] = 21'b100000000000000000000;
 buffer[1155] = 21'b100000000000000000000;
 buffer[1156] = 21'b100000000000000000000;
 buffer[1157] = 21'b100000000000000000000;
 buffer[1158] = 21'b100000000000000000000;
 buffer[1159] = 21'b100000000000000000000;
 buffer[1160] = 21'b100000000000000000000;
 buffer[1161] = 21'b100000000000000000000;
 buffer[1162] = 21'b100000000000000000000;
 buffer[1163] = 21'b100000000000000000000;
 buffer[1164] = 21'b100000000000000000000;
 buffer[1165] = 21'b100000000000000000000;
 buffer[1166] = 21'b100000000000000000000;
 buffer[1167] = 21'b100000000000000000000;
 buffer[1168] = 21'b100000000000000000000;
 buffer[1169] = 21'b100000000000000000000;
 buffer[1170] = 21'b100000000000000000000;
 buffer[1171] = 21'b100000000000000000000;
 buffer[1172] = 21'b100000000000000000000;
 buffer[1173] = 21'b100000000000000000000;
 buffer[1174] = 21'b100000000000000000000;
 buffer[1175] = 21'b100000000000000000000;
 buffer[1176] = 21'b100000000000000000000;
 buffer[1177] = 21'b100000000000000000000;
 buffer[1178] = 21'b100000000000000000000;
 buffer[1179] = 21'b100000000000000000000;
 buffer[1180] = 21'b100000000000000000000;
 buffer[1181] = 21'b100000000000000000000;
 buffer[1182] = 21'b100000000000000000000;
 buffer[1183] = 21'b100000000000000000000;
 buffer[1184] = 21'b100000000000000000000;
 buffer[1185] = 21'b100000000000000000000;
 buffer[1186] = 21'b100000000000000000000;
 buffer[1187] = 21'b100000000000000000000;
 buffer[1188] = 21'b100000000000000000000;
 buffer[1189] = 21'b100000000000000000000;
 buffer[1190] = 21'b100000000000000000000;
 buffer[1191] = 21'b100000000000000000000;
 buffer[1192] = 21'b100000000000000000000;
 buffer[1193] = 21'b100000000000000000000;
 buffer[1194] = 21'b100000000000000000000;
 buffer[1195] = 21'b100000000000000000000;
 buffer[1196] = 21'b100000000000000000000;
 buffer[1197] = 21'b100000000000000000000;
 buffer[1198] = 21'b100000000000000000000;
 buffer[1199] = 21'b100000000000000000000;
 buffer[1200] = 21'b100000000000000000000;
 buffer[1201] = 21'b100000000000000000000;
 buffer[1202] = 21'b100000000000000000000;
 buffer[1203] = 21'b100000000000000000000;
 buffer[1204] = 21'b100000000000000000000;
 buffer[1205] = 21'b100000000000000000000;
 buffer[1206] = 21'b100000000000000000000;
 buffer[1207] = 21'b100000000000000000000;
 buffer[1208] = 21'b100000000000000000000;
 buffer[1209] = 21'b100000000000000000000;
 buffer[1210] = 21'b100000000000000000000;
 buffer[1211] = 21'b100000000000000000000;
 buffer[1212] = 21'b100000000000000000000;
 buffer[1213] = 21'b100000000000000000000;
 buffer[1214] = 21'b100000000000000000000;
 buffer[1215] = 21'b100000000000000000000;
 buffer[1216] = 21'b100000000000000000000;
 buffer[1217] = 21'b100000000000000000000;
 buffer[1218] = 21'b100000000000000000000;
 buffer[1219] = 21'b100000000000000000000;
 buffer[1220] = 21'b100000000000000000000;
 buffer[1221] = 21'b100000000000000000000;
 buffer[1222] = 21'b100000000000000000000;
 buffer[1223] = 21'b100000000000000000000;
 buffer[1224] = 21'b100000000000000000000;
 buffer[1225] = 21'b100000000000000000000;
 buffer[1226] = 21'b100000000000000000000;
 buffer[1227] = 21'b100000000000000000000;
 buffer[1228] = 21'b100000000000000000000;
 buffer[1229] = 21'b100000000000000000000;
 buffer[1230] = 21'b100000000000000000000;
 buffer[1231] = 21'b100000000000000000000;
 buffer[1232] = 21'b100000000000000000000;
 buffer[1233] = 21'b100000000000000000000;
 buffer[1234] = 21'b100000000000000000000;
 buffer[1235] = 21'b100000000000000000000;
 buffer[1236] = 21'b100000000000000000000;
 buffer[1237] = 21'b100000000000000000000;
 buffer[1238] = 21'b100000000000000000000;
 buffer[1239] = 21'b100000000000000000000;
 buffer[1240] = 21'b100000000000000000000;
 buffer[1241] = 21'b100000000000000000000;
 buffer[1242] = 21'b100000000000000000000;
 buffer[1243] = 21'b100000000000000000000;
 buffer[1244] = 21'b100000000000000000000;
 buffer[1245] = 21'b100000000000000000000;
 buffer[1246] = 21'b100000000000000000000;
 buffer[1247] = 21'b100000000000000000000;
 buffer[1248] = 21'b100000000000000000000;
 buffer[1249] = 21'b100000000000000000000;
 buffer[1250] = 21'b100000000000000000000;
 buffer[1251] = 21'b100000000000000000000;
 buffer[1252] = 21'b100000000000000000000;
 buffer[1253] = 21'b100000000000000000000;
 buffer[1254] = 21'b100000000000000000000;
 buffer[1255] = 21'b100000000000000000000;
 buffer[1256] = 21'b100000000000000000000;
 buffer[1257] = 21'b100000000000000000000;
 buffer[1258] = 21'b100000000000000000000;
 buffer[1259] = 21'b100000000000000000000;
 buffer[1260] = 21'b100000000000000000000;
 buffer[1261] = 21'b100000000000000000000;
 buffer[1262] = 21'b100000000000000000000;
 buffer[1263] = 21'b100000000000000000000;
 buffer[1264] = 21'b100000000000000000000;
 buffer[1265] = 21'b100000000000000000000;
 buffer[1266] = 21'b100000000000000000000;
 buffer[1267] = 21'b100000000000000000000;
 buffer[1268] = 21'b100000000000000000000;
 buffer[1269] = 21'b100000000000000000000;
 buffer[1270] = 21'b100000000000000000000;
 buffer[1271] = 21'b100000000000000000000;
 buffer[1272] = 21'b100000000000000000000;
 buffer[1273] = 21'b100000000000000000000;
 buffer[1274] = 21'b100000000000000000000;
 buffer[1275] = 21'b100000000000000000000;
 buffer[1276] = 21'b100000000000000000000;
 buffer[1277] = 21'b100000000000000000000;
 buffer[1278] = 21'b100000000000000000000;
 buffer[1279] = 21'b100000000000000000000;
 buffer[1280] = 21'b100000000000000000000;
 buffer[1281] = 21'b100000000000000000000;
 buffer[1282] = 21'b100000000000000000000;
 buffer[1283] = 21'b100000000000000000000;
 buffer[1284] = 21'b100000000000000000000;
 buffer[1285] = 21'b100000000000000000000;
 buffer[1286] = 21'b100000000000000000000;
 buffer[1287] = 21'b100000000000000000000;
 buffer[1288] = 21'b100000000000000000000;
 buffer[1289] = 21'b100000000000000000000;
 buffer[1290] = 21'b100000000000000000000;
 buffer[1291] = 21'b100000000000000000000;
 buffer[1292] = 21'b100000000000000000000;
 buffer[1293] = 21'b100000000000000000000;
 buffer[1294] = 21'b100000000000000000000;
 buffer[1295] = 21'b100000000000000000000;
 buffer[1296] = 21'b100000000000000000000;
 buffer[1297] = 21'b100000000000000000000;
 buffer[1298] = 21'b100000000000000000000;
 buffer[1299] = 21'b100000000000000000000;
 buffer[1300] = 21'b100000000000000000000;
 buffer[1301] = 21'b100000000000000000000;
 buffer[1302] = 21'b100000000000000000000;
 buffer[1303] = 21'b100000000000000000000;
 buffer[1304] = 21'b100000000000000000000;
 buffer[1305] = 21'b100000000000000000000;
 buffer[1306] = 21'b100000000000000000000;
 buffer[1307] = 21'b100000000000000000000;
 buffer[1308] = 21'b100000000000000000000;
 buffer[1309] = 21'b100000000000000000000;
 buffer[1310] = 21'b100000000000000000000;
 buffer[1311] = 21'b100000000000000000000;
 buffer[1312] = 21'b100000000000000000000;
 buffer[1313] = 21'b100000000000000000000;
 buffer[1314] = 21'b100000000000000000000;
 buffer[1315] = 21'b100000000000000000000;
 buffer[1316] = 21'b100000000000000000000;
 buffer[1317] = 21'b100000000000000000000;
 buffer[1318] = 21'b100000000000000000000;
 buffer[1319] = 21'b100000000000000000000;
 buffer[1320] = 21'b100000000000000000000;
 buffer[1321] = 21'b100000000000000000000;
 buffer[1322] = 21'b100000000000000000000;
 buffer[1323] = 21'b100000000000000000000;
 buffer[1324] = 21'b100000000000000000000;
 buffer[1325] = 21'b100000000000000000000;
 buffer[1326] = 21'b100000000000000000000;
 buffer[1327] = 21'b100000000000000000000;
 buffer[1328] = 21'b100000000000000000000;
 buffer[1329] = 21'b100000000000000000000;
 buffer[1330] = 21'b100000000000000000000;
 buffer[1331] = 21'b100000000000000000000;
 buffer[1332] = 21'b100000000000000000000;
 buffer[1333] = 21'b100000000000000000000;
 buffer[1334] = 21'b100000000000000000000;
 buffer[1335] = 21'b100000000000000000000;
 buffer[1336] = 21'b100000000000000000000;
 buffer[1337] = 21'b100000000000000000000;
 buffer[1338] = 21'b100000000000000000000;
 buffer[1339] = 21'b100000000000000000000;
 buffer[1340] = 21'b100000000000000000000;
 buffer[1341] = 21'b100000000000000000000;
 buffer[1342] = 21'b100000000000000000000;
 buffer[1343] = 21'b100000000000000000000;
 buffer[1344] = 21'b100000000000000000000;
 buffer[1345] = 21'b100000000000000000000;
 buffer[1346] = 21'b100000000000000000000;
 buffer[1347] = 21'b100000000000000000000;
 buffer[1348] = 21'b100000000000000000000;
 buffer[1349] = 21'b100000000000000000000;
 buffer[1350] = 21'b100000000000000000000;
 buffer[1351] = 21'b100000000000000000000;
 buffer[1352] = 21'b100000000000000000000;
 buffer[1353] = 21'b100000000000000000000;
 buffer[1354] = 21'b100000000000000000000;
 buffer[1355] = 21'b100000000000000000000;
 buffer[1356] = 21'b100000000000000000000;
 buffer[1357] = 21'b100000000000000000000;
 buffer[1358] = 21'b100000000000000000000;
 buffer[1359] = 21'b100000000000000000000;
 buffer[1360] = 21'b100000000000000000000;
 buffer[1361] = 21'b100000000000000000000;
 buffer[1362] = 21'b100000000000000000000;
 buffer[1363] = 21'b100000000000000000000;
 buffer[1364] = 21'b100000000000000000000;
 buffer[1365] = 21'b100000000000000000000;
 buffer[1366] = 21'b100000000000000000000;
 buffer[1367] = 21'b100000000000000000000;
 buffer[1368] = 21'b100000000000000000000;
 buffer[1369] = 21'b100000000000000000000;
 buffer[1370] = 21'b100000000000000000000;
 buffer[1371] = 21'b100000000000000000000;
 buffer[1372] = 21'b100000000000000000000;
 buffer[1373] = 21'b100000000000000000000;
 buffer[1374] = 21'b100000000000000000000;
 buffer[1375] = 21'b100000000000000000000;
 buffer[1376] = 21'b100000000000000000000;
 buffer[1377] = 21'b100000000000000000000;
 buffer[1378] = 21'b100000000000000000000;
 buffer[1379] = 21'b100000000000000000000;
 buffer[1380] = 21'b100000000000000000000;
 buffer[1381] = 21'b100000000000000000000;
 buffer[1382] = 21'b100000000000000000000;
 buffer[1383] = 21'b100000000000000000000;
 buffer[1384] = 21'b100000000000000000000;
 buffer[1385] = 21'b100000000000000000000;
 buffer[1386] = 21'b100000000000000000000;
 buffer[1387] = 21'b100000000000000000000;
 buffer[1388] = 21'b100000000000000000000;
 buffer[1389] = 21'b100000000000000000000;
 buffer[1390] = 21'b100000000000000000000;
 buffer[1391] = 21'b100000000000000000000;
 buffer[1392] = 21'b100000000000000000000;
 buffer[1393] = 21'b100000000000000000000;
 buffer[1394] = 21'b100000000000000000000;
 buffer[1395] = 21'b100000000000000000000;
 buffer[1396] = 21'b100000000000000000000;
 buffer[1397] = 21'b100000000000000000000;
 buffer[1398] = 21'b100000000000000000000;
 buffer[1399] = 21'b100000000000000000000;
 buffer[1400] = 21'b100000000000000000000;
 buffer[1401] = 21'b100000000000000000000;
 buffer[1402] = 21'b100000000000000000000;
 buffer[1403] = 21'b100000000000000000000;
 buffer[1404] = 21'b100000000000000000000;
 buffer[1405] = 21'b100000000000000000000;
 buffer[1406] = 21'b100000000000000000000;
 buffer[1407] = 21'b100000000000000000000;
 buffer[1408] = 21'b100000000000000000000;
 buffer[1409] = 21'b100000000000000000000;
 buffer[1410] = 21'b100000000000000000000;
 buffer[1411] = 21'b100000000000000000000;
 buffer[1412] = 21'b100000000000000000000;
 buffer[1413] = 21'b100000000000000000000;
 buffer[1414] = 21'b100000000000000000000;
 buffer[1415] = 21'b100000000000000000000;
 buffer[1416] = 21'b100000000000000000000;
 buffer[1417] = 21'b100000000000000000000;
 buffer[1418] = 21'b100000000000000000000;
 buffer[1419] = 21'b100000000000000000000;
 buffer[1420] = 21'b100000000000000000000;
 buffer[1421] = 21'b100000000000000000000;
 buffer[1422] = 21'b100000000000000000000;
 buffer[1423] = 21'b100000000000000000000;
 buffer[1424] = 21'b100000000000000000000;
 buffer[1425] = 21'b100000000000000000000;
 buffer[1426] = 21'b100000000000000000000;
 buffer[1427] = 21'b100000000000000000000;
 buffer[1428] = 21'b100000000000000000000;
 buffer[1429] = 21'b100000000000000000000;
 buffer[1430] = 21'b100000000000000000000;
 buffer[1431] = 21'b100000000000000000000;
 buffer[1432] = 21'b100000000000000000000;
 buffer[1433] = 21'b100000000000000000000;
 buffer[1434] = 21'b100000000000000000000;
 buffer[1435] = 21'b100000000000000000000;
 buffer[1436] = 21'b100000000000000000000;
 buffer[1437] = 21'b100000000000000000000;
 buffer[1438] = 21'b100000000000000000000;
 buffer[1439] = 21'b100000000000000000000;
 buffer[1440] = 21'b100000000000000000000;
 buffer[1441] = 21'b100000000000000000000;
 buffer[1442] = 21'b100000000000000000000;
 buffer[1443] = 21'b100000000000000000000;
 buffer[1444] = 21'b100000000000000000000;
 buffer[1445] = 21'b100000000000000000000;
 buffer[1446] = 21'b100000000000000000000;
 buffer[1447] = 21'b100000000000000000000;
 buffer[1448] = 21'b100000000000000000000;
 buffer[1449] = 21'b100000000000000000000;
 buffer[1450] = 21'b100000000000000000000;
 buffer[1451] = 21'b100000000000000000000;
 buffer[1452] = 21'b100000000000000000000;
 buffer[1453] = 21'b100000000000000000000;
 buffer[1454] = 21'b100000000000000000000;
 buffer[1455] = 21'b100000000000000000000;
 buffer[1456] = 21'b100000000000000000000;
 buffer[1457] = 21'b100000000000000000000;
 buffer[1458] = 21'b100000000000000000000;
 buffer[1459] = 21'b100000000000000000000;
 buffer[1460] = 21'b100000000000000000000;
 buffer[1461] = 21'b100000000000000000000;
 buffer[1462] = 21'b100000000000000000000;
 buffer[1463] = 21'b100000000000000000000;
 buffer[1464] = 21'b100000000000000000000;
 buffer[1465] = 21'b100000000000000000000;
 buffer[1466] = 21'b100000000000000000000;
 buffer[1467] = 21'b100000000000000000000;
 buffer[1468] = 21'b100000000000000000000;
 buffer[1469] = 21'b100000000000000000000;
 buffer[1470] = 21'b100000000000000000000;
 buffer[1471] = 21'b100000000000000000000;
 buffer[1472] = 21'b100000000000000000000;
 buffer[1473] = 21'b100000000000000000000;
 buffer[1474] = 21'b100000000000000000000;
 buffer[1475] = 21'b100000000000000000000;
 buffer[1476] = 21'b100000000000000000000;
 buffer[1477] = 21'b100000000000000000000;
 buffer[1478] = 21'b100000000000000000000;
 buffer[1479] = 21'b100000000000000000000;
 buffer[1480] = 21'b100000000000000000000;
 buffer[1481] = 21'b100000000000000000000;
 buffer[1482] = 21'b100000000000000000000;
 buffer[1483] = 21'b100000000000000000000;
 buffer[1484] = 21'b100000000000000000000;
 buffer[1485] = 21'b100000000000000000000;
 buffer[1486] = 21'b100000000000000000000;
 buffer[1487] = 21'b100000000000000000000;
 buffer[1488] = 21'b100000000000000000000;
 buffer[1489] = 21'b100000000000000000000;
 buffer[1490] = 21'b100000000000000000000;
 buffer[1491] = 21'b100000000000000000000;
 buffer[1492] = 21'b100000000000000000000;
 buffer[1493] = 21'b100000000000000000000;
 buffer[1494] = 21'b100000000000000000000;
 buffer[1495] = 21'b100000000000000000000;
 buffer[1496] = 21'b100000000000000000000;
 buffer[1497] = 21'b100000000000000000000;
 buffer[1498] = 21'b100000000000000000000;
 buffer[1499] = 21'b100000000000000000000;
 buffer[1500] = 21'b100000000000000000000;
 buffer[1501] = 21'b100000000000000000000;
 buffer[1502] = 21'b100000000000000000000;
 buffer[1503] = 21'b100000000000000000000;
 buffer[1504] = 21'b100000000000000000000;
 buffer[1505] = 21'b100000000000000000000;
 buffer[1506] = 21'b100000000000000000000;
 buffer[1507] = 21'b100000000000000000000;
 buffer[1508] = 21'b100000000000000000000;
 buffer[1509] = 21'b100000000000000000000;
 buffer[1510] = 21'b100000000000000000000;
 buffer[1511] = 21'b100000000000000000000;
 buffer[1512] = 21'b100000000000000000000;
 buffer[1513] = 21'b100000000000000000000;
 buffer[1514] = 21'b100000000000000000000;
 buffer[1515] = 21'b100000000000000000000;
 buffer[1516] = 21'b100000000000000000000;
 buffer[1517] = 21'b100000000000000000000;
 buffer[1518] = 21'b100000000000000000000;
 buffer[1519] = 21'b100000000000000000000;
 buffer[1520] = 21'b100000000000000000000;
 buffer[1521] = 21'b100000000000000000000;
 buffer[1522] = 21'b100000000000000000000;
 buffer[1523] = 21'b100000000000000000000;
 buffer[1524] = 21'b100000000000000000000;
 buffer[1525] = 21'b100000000000000000000;
 buffer[1526] = 21'b100000000000000000000;
 buffer[1527] = 21'b100000000000000000000;
 buffer[1528] = 21'b100000000000000000000;
 buffer[1529] = 21'b100000000000000000000;
 buffer[1530] = 21'b100000000000000000000;
 buffer[1531] = 21'b100000000000000000000;
 buffer[1532] = 21'b100000000000000000000;
 buffer[1533] = 21'b100000000000000000000;
 buffer[1534] = 21'b100000000000000000000;
 buffer[1535] = 21'b100000000000000000000;
 buffer[1536] = 21'b100000000000000000000;
 buffer[1537] = 21'b100000000000000000000;
 buffer[1538] = 21'b100000000000000000000;
 buffer[1539] = 21'b100000000000000000000;
 buffer[1540] = 21'b100000000000000000000;
 buffer[1541] = 21'b100000000000000000000;
 buffer[1542] = 21'b100000000000000000000;
 buffer[1543] = 21'b100000000000000000000;
 buffer[1544] = 21'b100000000000000000000;
 buffer[1545] = 21'b100000000000000000000;
 buffer[1546] = 21'b100000000000000000000;
 buffer[1547] = 21'b100000000000000000000;
 buffer[1548] = 21'b100000000000000000000;
 buffer[1549] = 21'b100000000000000000000;
 buffer[1550] = 21'b100000000000000000000;
 buffer[1551] = 21'b100000000000000000000;
 buffer[1552] = 21'b100000000000000000000;
 buffer[1553] = 21'b100000000000000000000;
 buffer[1554] = 21'b100000000000000000000;
 buffer[1555] = 21'b100000000000000000000;
 buffer[1556] = 21'b100000000000000000000;
 buffer[1557] = 21'b100000000000000000000;
 buffer[1558] = 21'b100000000000000000000;
 buffer[1559] = 21'b100000000000000000000;
 buffer[1560] = 21'b100000000000000000000;
 buffer[1561] = 21'b100000000000000000000;
 buffer[1562] = 21'b100000000000000000000;
 buffer[1563] = 21'b100000000000000000000;
 buffer[1564] = 21'b100000000000000000000;
 buffer[1565] = 21'b100000000000000000000;
 buffer[1566] = 21'b100000000000000000000;
 buffer[1567] = 21'b100000000000000000000;
 buffer[1568] = 21'b100000000000000000000;
 buffer[1569] = 21'b100000000000000000000;
 buffer[1570] = 21'b100000000000000000000;
 buffer[1571] = 21'b100000000000000000000;
 buffer[1572] = 21'b100000000000000000000;
 buffer[1573] = 21'b100000000000000000000;
 buffer[1574] = 21'b100000000000000000000;
 buffer[1575] = 21'b100000000000000000000;
 buffer[1576] = 21'b100000000000000000000;
 buffer[1577] = 21'b100000000000000000000;
 buffer[1578] = 21'b100000000000000000000;
 buffer[1579] = 21'b100000000000000000000;
 buffer[1580] = 21'b100000000000000000000;
 buffer[1581] = 21'b100000000000000000000;
 buffer[1582] = 21'b100000000000000000000;
 buffer[1583] = 21'b100000000000000000000;
 buffer[1584] = 21'b100000000000000000000;
 buffer[1585] = 21'b100000000000000000000;
 buffer[1586] = 21'b100000000000000000000;
 buffer[1587] = 21'b100000000000000000000;
 buffer[1588] = 21'b100000000000000000000;
 buffer[1589] = 21'b100000000000000000000;
 buffer[1590] = 21'b100000000000000000000;
 buffer[1591] = 21'b100000000000000000000;
 buffer[1592] = 21'b100000000000000000000;
 buffer[1593] = 21'b100000000000000000000;
 buffer[1594] = 21'b100000000000000000000;
 buffer[1595] = 21'b100000000000000000000;
 buffer[1596] = 21'b100000000000000000000;
 buffer[1597] = 21'b100000000000000000000;
 buffer[1598] = 21'b100000000000000000000;
 buffer[1599] = 21'b100000000000000000000;
 buffer[1600] = 21'b100000000000000000000;
 buffer[1601] = 21'b100000000000000000000;
 buffer[1602] = 21'b100000000000000000000;
 buffer[1603] = 21'b100000000000000000000;
 buffer[1604] = 21'b100000000000000000000;
 buffer[1605] = 21'b100000000000000000000;
 buffer[1606] = 21'b100000000000000000000;
 buffer[1607] = 21'b100000000000000000000;
 buffer[1608] = 21'b100000000000000000000;
 buffer[1609] = 21'b100000000000000000000;
 buffer[1610] = 21'b100000000000000000000;
 buffer[1611] = 21'b100000000000000000000;
 buffer[1612] = 21'b100000000000000000000;
 buffer[1613] = 21'b100000000000000000000;
 buffer[1614] = 21'b100000000000000000000;
 buffer[1615] = 21'b100000000000000000000;
 buffer[1616] = 21'b100000000000000000000;
 buffer[1617] = 21'b100000000000000000000;
 buffer[1618] = 21'b100000000000000000000;
 buffer[1619] = 21'b100000000000000000000;
 buffer[1620] = 21'b100000000000000000000;
 buffer[1621] = 21'b100000000000000000000;
 buffer[1622] = 21'b100000000000000000000;
 buffer[1623] = 21'b100000000000000000000;
 buffer[1624] = 21'b100000000000000000000;
 buffer[1625] = 21'b100000000000000000000;
 buffer[1626] = 21'b100000000000000000000;
 buffer[1627] = 21'b100000000000000000000;
 buffer[1628] = 21'b100000000000000000000;
 buffer[1629] = 21'b100000000000000000000;
 buffer[1630] = 21'b100000000000000000000;
 buffer[1631] = 21'b100000000000000000000;
 buffer[1632] = 21'b100000000000000000000;
 buffer[1633] = 21'b100000000000000000000;
 buffer[1634] = 21'b100000000000000000000;
 buffer[1635] = 21'b100000000000000000000;
 buffer[1636] = 21'b100000000000000000000;
 buffer[1637] = 21'b100000000000000000000;
 buffer[1638] = 21'b100000000000000000000;
 buffer[1639] = 21'b100000000000000000000;
 buffer[1640] = 21'b100000000000000000000;
 buffer[1641] = 21'b100000000000000000000;
 buffer[1642] = 21'b100000000000000000000;
 buffer[1643] = 21'b100000000000000000000;
 buffer[1644] = 21'b100000000000000000000;
 buffer[1645] = 21'b100000000000000000000;
 buffer[1646] = 21'b100000000000000000000;
 buffer[1647] = 21'b100000000000000000000;
 buffer[1648] = 21'b100000000000000000000;
 buffer[1649] = 21'b100000000000000000000;
 buffer[1650] = 21'b100000000000000000000;
 buffer[1651] = 21'b100000000000000000000;
 buffer[1652] = 21'b100000000000000000000;
 buffer[1653] = 21'b100000000000000000000;
 buffer[1654] = 21'b100000000000000000000;
 buffer[1655] = 21'b100000000000000000000;
 buffer[1656] = 21'b100000000000000000000;
 buffer[1657] = 21'b100000000000000000000;
 buffer[1658] = 21'b100000000000000000000;
 buffer[1659] = 21'b100000000000000000000;
 buffer[1660] = 21'b100000000000000000000;
 buffer[1661] = 21'b100000000000000000000;
 buffer[1662] = 21'b100000000000000000000;
 buffer[1663] = 21'b100000000000000000000;
 buffer[1664] = 21'b100000000000000000000;
 buffer[1665] = 21'b100000000000000000000;
 buffer[1666] = 21'b100000000000000000000;
 buffer[1667] = 21'b100000000000000000000;
 buffer[1668] = 21'b100000000000000000000;
 buffer[1669] = 21'b100000000000000000000;
 buffer[1670] = 21'b100000000000000000000;
 buffer[1671] = 21'b100000000000000000000;
 buffer[1672] = 21'b100000000000000000000;
 buffer[1673] = 21'b100000000000000000000;
 buffer[1674] = 21'b100000000000000000000;
 buffer[1675] = 21'b100000000000000000000;
 buffer[1676] = 21'b100000000000000000000;
 buffer[1677] = 21'b100000000000000000000;
 buffer[1678] = 21'b100000000000000000000;
 buffer[1679] = 21'b100000000000000000000;
 buffer[1680] = 21'b100000000000000000000;
 buffer[1681] = 21'b100000000000000000000;
 buffer[1682] = 21'b100000000000000000000;
 buffer[1683] = 21'b100000000000000000000;
 buffer[1684] = 21'b100000000000000000000;
 buffer[1685] = 21'b100000000000000000000;
 buffer[1686] = 21'b100000000000000000000;
 buffer[1687] = 21'b100000000000000000000;
 buffer[1688] = 21'b100000000000000000000;
 buffer[1689] = 21'b100000000000000000000;
 buffer[1690] = 21'b100000000000000000000;
 buffer[1691] = 21'b100000000000000000000;
 buffer[1692] = 21'b100000000000000000000;
 buffer[1693] = 21'b100000000000000000000;
 buffer[1694] = 21'b100000000000000000000;
 buffer[1695] = 21'b100000000000000000000;
 buffer[1696] = 21'b100000000000000000000;
 buffer[1697] = 21'b100000000000000000000;
 buffer[1698] = 21'b100000000000000000000;
 buffer[1699] = 21'b100000000000000000000;
 buffer[1700] = 21'b100000000000000000000;
 buffer[1701] = 21'b100000000000000000000;
 buffer[1702] = 21'b100000000000000000000;
 buffer[1703] = 21'b100000000000000000000;
 buffer[1704] = 21'b100000000000000000000;
 buffer[1705] = 21'b100000000000000000000;
 buffer[1706] = 21'b100000000000000000000;
 buffer[1707] = 21'b100000000000000000000;
 buffer[1708] = 21'b100000000000000000000;
 buffer[1709] = 21'b100000000000000000000;
 buffer[1710] = 21'b100000000000000000000;
 buffer[1711] = 21'b100000000000000000000;
 buffer[1712] = 21'b100000000000000000000;
 buffer[1713] = 21'b100000000000000000000;
 buffer[1714] = 21'b100000000000000000000;
 buffer[1715] = 21'b100000000000000000000;
 buffer[1716] = 21'b100000000000000000000;
 buffer[1717] = 21'b100000000000000000000;
 buffer[1718] = 21'b100000000000000000000;
 buffer[1719] = 21'b100000000000000000000;
 buffer[1720] = 21'b100000000000000000000;
 buffer[1721] = 21'b100000000000000000000;
 buffer[1722] = 21'b100000000000000000000;
 buffer[1723] = 21'b100000000000000000000;
 buffer[1724] = 21'b100000000000000000000;
 buffer[1725] = 21'b100000000000000000000;
 buffer[1726] = 21'b100000000000000000000;
 buffer[1727] = 21'b100000000000000000000;
 buffer[1728] = 21'b100000000000000000000;
 buffer[1729] = 21'b100000000000000000000;
 buffer[1730] = 21'b100000000000000000000;
 buffer[1731] = 21'b100000000000000000000;
 buffer[1732] = 21'b100000000000000000000;
 buffer[1733] = 21'b100000000000000000000;
 buffer[1734] = 21'b100000000000000000000;
 buffer[1735] = 21'b100000000000000000000;
 buffer[1736] = 21'b100000000000000000000;
 buffer[1737] = 21'b100000000000000000000;
 buffer[1738] = 21'b100000000000000000000;
 buffer[1739] = 21'b100000000000000000000;
 buffer[1740] = 21'b100000000000000000000;
 buffer[1741] = 21'b100000000000000000000;
 buffer[1742] = 21'b100000000000000000000;
 buffer[1743] = 21'b100000000000000000000;
 buffer[1744] = 21'b100000000000000000000;
 buffer[1745] = 21'b100000000000000000000;
 buffer[1746] = 21'b100000000000000000000;
 buffer[1747] = 21'b100000000000000000000;
 buffer[1748] = 21'b100000000000000000000;
 buffer[1749] = 21'b100000000000000000000;
 buffer[1750] = 21'b100000000000000000000;
 buffer[1751] = 21'b100000000000000000000;
 buffer[1752] = 21'b100000000000000000000;
 buffer[1753] = 21'b100000000000000000000;
 buffer[1754] = 21'b100000000000000000000;
 buffer[1755] = 21'b100000000000000000000;
 buffer[1756] = 21'b100000000000000000000;
 buffer[1757] = 21'b100000000000000000000;
 buffer[1758] = 21'b100000000000000000000;
 buffer[1759] = 21'b100000000000000000000;
 buffer[1760] = 21'b100000000000000000000;
 buffer[1761] = 21'b100000000000000000000;
 buffer[1762] = 21'b100000000000000000000;
 buffer[1763] = 21'b100000000000000000000;
 buffer[1764] = 21'b100000000000000000000;
 buffer[1765] = 21'b100000000000000000000;
 buffer[1766] = 21'b100000000000000000000;
 buffer[1767] = 21'b100000000000000000000;
 buffer[1768] = 21'b100000000000000000000;
 buffer[1769] = 21'b100000000000000000000;
 buffer[1770] = 21'b100000000000000000000;
 buffer[1771] = 21'b100000000000000000000;
 buffer[1772] = 21'b100000000000000000000;
 buffer[1773] = 21'b100000000000000000000;
 buffer[1774] = 21'b100000000000000000000;
 buffer[1775] = 21'b100000000000000000000;
 buffer[1776] = 21'b100000000000000000000;
 buffer[1777] = 21'b100000000000000000000;
 buffer[1778] = 21'b100000000000000000000;
 buffer[1779] = 21'b100000000000000000000;
 buffer[1780] = 21'b100000000000000000000;
 buffer[1781] = 21'b100000000000000000000;
 buffer[1782] = 21'b100000000000000000000;
 buffer[1783] = 21'b100000000000000000000;
 buffer[1784] = 21'b100000000000000000000;
 buffer[1785] = 21'b100000000000000000000;
 buffer[1786] = 21'b100000000000000000000;
 buffer[1787] = 21'b100000000000000000000;
 buffer[1788] = 21'b100000000000000000000;
 buffer[1789] = 21'b100000000000000000000;
 buffer[1790] = 21'b100000000000000000000;
 buffer[1791] = 21'b100000000000000000000;
 buffer[1792] = 21'b100000000000000000000;
 buffer[1793] = 21'b100000000000000000000;
 buffer[1794] = 21'b100000000000000000000;
 buffer[1795] = 21'b100000000000000000000;
 buffer[1796] = 21'b100000000000000000000;
 buffer[1797] = 21'b100000000000000000000;
 buffer[1798] = 21'b100000000000000000000;
 buffer[1799] = 21'b100000000000000000000;
 buffer[1800] = 21'b100000000000000000000;
 buffer[1801] = 21'b100000000000000000000;
 buffer[1802] = 21'b100000000000000000000;
 buffer[1803] = 21'b100000000000000000000;
 buffer[1804] = 21'b100000000000000000000;
 buffer[1805] = 21'b100000000000000000000;
 buffer[1806] = 21'b100000000000000000000;
 buffer[1807] = 21'b100000000000000000000;
 buffer[1808] = 21'b100000000000000000000;
 buffer[1809] = 21'b100000000000000000000;
 buffer[1810] = 21'b100000000000000000000;
 buffer[1811] = 21'b100000000000000000000;
 buffer[1812] = 21'b100000000000000000000;
 buffer[1813] = 21'b100000000000000000000;
 buffer[1814] = 21'b100000000000000000000;
 buffer[1815] = 21'b100000000000000000000;
 buffer[1816] = 21'b100000000000000000000;
 buffer[1817] = 21'b100000000000000000000;
 buffer[1818] = 21'b100000000000000000000;
 buffer[1819] = 21'b100000000000000000000;
 buffer[1820] = 21'b100000000000000000000;
 buffer[1821] = 21'b100000000000000000000;
 buffer[1822] = 21'b100000000000000000000;
 buffer[1823] = 21'b100000000000000000000;
 buffer[1824] = 21'b100000000000000000000;
 buffer[1825] = 21'b100000000000000000000;
 buffer[1826] = 21'b100000000000000000000;
 buffer[1827] = 21'b100000000000000000000;
 buffer[1828] = 21'b100000000000000000000;
 buffer[1829] = 21'b100000000000000000000;
 buffer[1830] = 21'b100000000000000000000;
 buffer[1831] = 21'b100000000000000000000;
 buffer[1832] = 21'b100000000000000000000;
 buffer[1833] = 21'b100000000000000000000;
 buffer[1834] = 21'b100000000000000000000;
 buffer[1835] = 21'b100000000000000000000;
 buffer[1836] = 21'b100000000000000000000;
 buffer[1837] = 21'b100000000000000000000;
 buffer[1838] = 21'b100000000000000000000;
 buffer[1839] = 21'b100000000000000000000;
 buffer[1840] = 21'b100000000000000000000;
 buffer[1841] = 21'b100000000000000000000;
 buffer[1842] = 21'b100000000000000000000;
 buffer[1843] = 21'b100000000000000000000;
 buffer[1844] = 21'b100000000000000000000;
 buffer[1845] = 21'b100000000000000000000;
 buffer[1846] = 21'b100000000000000000000;
 buffer[1847] = 21'b100000000000000000000;
 buffer[1848] = 21'b100000000000000000000;
 buffer[1849] = 21'b100000000000000000000;
 buffer[1850] = 21'b100000000000000000000;
 buffer[1851] = 21'b100000000000000000000;
 buffer[1852] = 21'b100000000000000000000;
 buffer[1853] = 21'b100000000000000000000;
 buffer[1854] = 21'b100000000000000000000;
 buffer[1855] = 21'b100000000000000000000;
 buffer[1856] = 21'b100000000000000000000;
 buffer[1857] = 21'b100000000000000000000;
 buffer[1858] = 21'b100000000000000000000;
 buffer[1859] = 21'b100000000000000000000;
 buffer[1860] = 21'b100000000000000000000;
 buffer[1861] = 21'b100000000000000000000;
 buffer[1862] = 21'b100000000000000000000;
 buffer[1863] = 21'b100000000000000000000;
 buffer[1864] = 21'b100000000000000000000;
 buffer[1865] = 21'b100000000000000000000;
 buffer[1866] = 21'b100000000000000000000;
 buffer[1867] = 21'b100000000000000000000;
 buffer[1868] = 21'b100000000000000000000;
 buffer[1869] = 21'b100000000000000000000;
 buffer[1870] = 21'b100000000000000000000;
 buffer[1871] = 21'b100000000000000000000;
 buffer[1872] = 21'b100000000000000000000;
 buffer[1873] = 21'b100000000000000000000;
 buffer[1874] = 21'b100000000000000000000;
 buffer[1875] = 21'b100000000000000000000;
 buffer[1876] = 21'b100000000000000000000;
 buffer[1877] = 21'b100000000000000000000;
 buffer[1878] = 21'b100000000000000000000;
 buffer[1879] = 21'b100000000000000000000;
 buffer[1880] = 21'b100000000000000000000;
 buffer[1881] = 21'b100000000000000000000;
 buffer[1882] = 21'b100000000000000000000;
 buffer[1883] = 21'b100000000000000000000;
 buffer[1884] = 21'b100000000000000000000;
 buffer[1885] = 21'b100000000000000000000;
 buffer[1886] = 21'b100000000000000000000;
 buffer[1887] = 21'b100000000000000000000;
 buffer[1888] = 21'b100000000000000000000;
 buffer[1889] = 21'b100000000000000000000;
 buffer[1890] = 21'b100000000000000000000;
 buffer[1891] = 21'b100000000000000000000;
 buffer[1892] = 21'b100000000000000000000;
 buffer[1893] = 21'b100000000000000000000;
 buffer[1894] = 21'b100000000000000000000;
 buffer[1895] = 21'b100000000000000000000;
 buffer[1896] = 21'b100000000000000000000;
 buffer[1897] = 21'b100000000000000000000;
 buffer[1898] = 21'b100000000000000000000;
 buffer[1899] = 21'b100000000000000000000;
 buffer[1900] = 21'b100000000000000000000;
 buffer[1901] = 21'b100000000000000000000;
 buffer[1902] = 21'b100000000000000000000;
 buffer[1903] = 21'b100000000000000000000;
 buffer[1904] = 21'b100000000000000000000;
 buffer[1905] = 21'b100000000000000000000;
 buffer[1906] = 21'b100000000000000000000;
 buffer[1907] = 21'b100000000000000000000;
 buffer[1908] = 21'b100000000000000000000;
 buffer[1909] = 21'b100000000000000000000;
 buffer[1910] = 21'b100000000000000000000;
 buffer[1911] = 21'b100000000000000000000;
 buffer[1912] = 21'b100000000000000000000;
 buffer[1913] = 21'b100000000000000000000;
 buffer[1914] = 21'b100000000000000000000;
 buffer[1915] = 21'b100000000000000000000;
 buffer[1916] = 21'b100000000000000000000;
 buffer[1917] = 21'b100000000000000000000;
 buffer[1918] = 21'b100000000000000000000;
 buffer[1919] = 21'b100000000000000000000;
 buffer[1920] = 21'b100000000000000000000;
 buffer[1921] = 21'b100000000000000000000;
 buffer[1922] = 21'b100000000000000000000;
 buffer[1923] = 21'b100000000000000000000;
 buffer[1924] = 21'b100000000000000000000;
 buffer[1925] = 21'b100000000000000000000;
 buffer[1926] = 21'b100000000000000000000;
 buffer[1927] = 21'b100000000000000000000;
 buffer[1928] = 21'b100000000000000000000;
 buffer[1929] = 21'b100000000000000000000;
 buffer[1930] = 21'b100000000000000000000;
 buffer[1931] = 21'b100000000000000000000;
 buffer[1932] = 21'b100000000000000000000;
 buffer[1933] = 21'b100000000000000000000;
 buffer[1934] = 21'b100000000000000000000;
 buffer[1935] = 21'b100000000000000000000;
 buffer[1936] = 21'b100000000000000000000;
 buffer[1937] = 21'b100000000000000000000;
 buffer[1938] = 21'b100000000000000000000;
 buffer[1939] = 21'b100000000000000000000;
 buffer[1940] = 21'b100000000000000000000;
 buffer[1941] = 21'b100000000000000000000;
 buffer[1942] = 21'b100000000000000000000;
 buffer[1943] = 21'b100000000000000000000;
 buffer[1944] = 21'b100000000000000000000;
 buffer[1945] = 21'b100000000000000000000;
 buffer[1946] = 21'b100000000000000000000;
 buffer[1947] = 21'b100000000000000000000;
 buffer[1948] = 21'b100000000000000000000;
 buffer[1949] = 21'b100000000000000000000;
 buffer[1950] = 21'b100000000000000000000;
 buffer[1951] = 21'b100000000000000000000;
 buffer[1952] = 21'b100000000000000000000;
 buffer[1953] = 21'b100000000000000000000;
 buffer[1954] = 21'b100000000000000000000;
 buffer[1955] = 21'b100000000000000000000;
 buffer[1956] = 21'b100000000000000000000;
 buffer[1957] = 21'b100000000000000000000;
 buffer[1958] = 21'b100000000000000000000;
 buffer[1959] = 21'b100000000000000000000;
 buffer[1960] = 21'b100000000000000000000;
 buffer[1961] = 21'b100000000000000000000;
 buffer[1962] = 21'b100000000000000000000;
 buffer[1963] = 21'b100000000000000000000;
 buffer[1964] = 21'b100000000000000000000;
 buffer[1965] = 21'b100000000000000000000;
 buffer[1966] = 21'b100000000000000000000;
 buffer[1967] = 21'b100000000000000000000;
 buffer[1968] = 21'b100000000000000000000;
 buffer[1969] = 21'b100000000000000000000;
 buffer[1970] = 21'b100000000000000000000;
 buffer[1971] = 21'b100000000000000000000;
 buffer[1972] = 21'b100000000000000000000;
 buffer[1973] = 21'b100000000000000000000;
 buffer[1974] = 21'b100000000000000000000;
 buffer[1975] = 21'b100000000000000000000;
 buffer[1976] = 21'b100000000000000000000;
 buffer[1977] = 21'b100000000000000000000;
 buffer[1978] = 21'b100000000000000000000;
 buffer[1979] = 21'b100000000000000000000;
 buffer[1980] = 21'b100000000000000000000;
 buffer[1981] = 21'b100000000000000000000;
 buffer[1982] = 21'b100000000000000000000;
 buffer[1983] = 21'b100000000000000000000;
 buffer[1984] = 21'b100000000000000000000;
 buffer[1985] = 21'b100000000000000000000;
 buffer[1986] = 21'b100000000000000000000;
 buffer[1987] = 21'b100000000000000000000;
 buffer[1988] = 21'b100000000000000000000;
 buffer[1989] = 21'b100000000000000000000;
 buffer[1990] = 21'b100000000000000000000;
 buffer[1991] = 21'b100000000000000000000;
 buffer[1992] = 21'b100000000000000000000;
 buffer[1993] = 21'b100000000000000000000;
 buffer[1994] = 21'b100000000000000000000;
 buffer[1995] = 21'b100000000000000000000;
 buffer[1996] = 21'b100000000000000000000;
 buffer[1997] = 21'b100000000000000000000;
 buffer[1998] = 21'b100000000000000000000;
 buffer[1999] = 21'b100000000000000000000;
 buffer[2000] = 21'b100000000000000000000;
 buffer[2001] = 21'b100000000000000000000;
 buffer[2002] = 21'b100000000000000000000;
 buffer[2003] = 21'b100000000000000000000;
 buffer[2004] = 21'b100000000000000000000;
 buffer[2005] = 21'b100000000000000000000;
 buffer[2006] = 21'b100000000000000000000;
 buffer[2007] = 21'b100000000000000000000;
 buffer[2008] = 21'b100000000000000000000;
 buffer[2009] = 21'b100000000000000000000;
 buffer[2010] = 21'b100000000000000000000;
 buffer[2011] = 21'b100000000000000000000;
 buffer[2012] = 21'b100000000000000000000;
 buffer[2013] = 21'b100000000000000000000;
 buffer[2014] = 21'b100000000000000000000;
 buffer[2015] = 21'b100000000000000000000;
 buffer[2016] = 21'b100000000000000000000;
 buffer[2017] = 21'b100000000000000000000;
 buffer[2018] = 21'b100000000000000000000;
 buffer[2019] = 21'b100000000000000000000;
 buffer[2020] = 21'b100000000000000000000;
 buffer[2021] = 21'b100000000000000000000;
 buffer[2022] = 21'b100000000000000000000;
 buffer[2023] = 21'b100000000000000000000;
 buffer[2024] = 21'b100000000000000000000;
 buffer[2025] = 21'b100000000000000000000;
 buffer[2026] = 21'b100000000000000000000;
 buffer[2027] = 21'b100000000000000000000;
 buffer[2028] = 21'b100000000000000000000;
 buffer[2029] = 21'b100000000000000000000;
 buffer[2030] = 21'b100000000000000000000;
 buffer[2031] = 21'b100000000000000000000;
 buffer[2032] = 21'b100000000000000000000;
 buffer[2033] = 21'b100000000000000000000;
 buffer[2034] = 21'b100000000000000000000;
 buffer[2035] = 21'b100000000000000000000;
 buffer[2036] = 21'b100000000000000000000;
 buffer[2037] = 21'b100000000000000000000;
 buffer[2038] = 21'b100000000000000000000;
 buffer[2039] = 21'b100000000000000000000;
 buffer[2040] = 21'b100000000000000000000;
 buffer[2041] = 21'b100000000000000000000;
 buffer[2042] = 21'b100000000000000000000;
 buffer[2043] = 21'b100000000000000000000;
 buffer[2044] = 21'b100000000000000000000;
 buffer[2045] = 21'b100000000000000000000;
 buffer[2046] = 21'b100000000000000000000;
 buffer[2047] = 21'b100000000000000000000;
 buffer[2048] = 21'b100000000000000000000;
 buffer[2049] = 21'b100000000000000000000;
 buffer[2050] = 21'b100000000000000000000;
 buffer[2051] = 21'b100000000000000000000;
 buffer[2052] = 21'b100000000000000000000;
 buffer[2053] = 21'b100000000000000000000;
 buffer[2054] = 21'b100000000000000000000;
 buffer[2055] = 21'b100000000000000000000;
 buffer[2056] = 21'b100000000000000000000;
 buffer[2057] = 21'b100000000000000000000;
 buffer[2058] = 21'b100000000000000000000;
 buffer[2059] = 21'b100000000000000000000;
 buffer[2060] = 21'b100000000000000000000;
 buffer[2061] = 21'b100000000000000000000;
 buffer[2062] = 21'b100000000000000000000;
 buffer[2063] = 21'b100000000000000000000;
 buffer[2064] = 21'b100000000000000000000;
 buffer[2065] = 21'b100000000000000000000;
 buffer[2066] = 21'b100000000000000000000;
 buffer[2067] = 21'b100000000000000000000;
 buffer[2068] = 21'b100000000000000000000;
 buffer[2069] = 21'b100000000000000000000;
 buffer[2070] = 21'b100000000000000000000;
 buffer[2071] = 21'b100000000000000000000;
 buffer[2072] = 21'b100000000000000000000;
 buffer[2073] = 21'b100000000000000000000;
 buffer[2074] = 21'b100000000000000000000;
 buffer[2075] = 21'b100000000000000000000;
 buffer[2076] = 21'b100000000000000000000;
 buffer[2077] = 21'b100000000000000000000;
 buffer[2078] = 21'b100000000000000000000;
 buffer[2079] = 21'b100000000000000000000;
 buffer[2080] = 21'b100000000000000000000;
 buffer[2081] = 21'b100000000000000000000;
 buffer[2082] = 21'b100000000000000000000;
 buffer[2083] = 21'b100000000000000000000;
 buffer[2084] = 21'b100000000000000000000;
 buffer[2085] = 21'b100000000000000000000;
 buffer[2086] = 21'b100000000000000000000;
 buffer[2087] = 21'b100000000000000000000;
 buffer[2088] = 21'b100000000000000000000;
 buffer[2089] = 21'b100000000000000000000;
 buffer[2090] = 21'b100000000000000000000;
 buffer[2091] = 21'b100000000000000000000;
 buffer[2092] = 21'b100000000000000000000;
 buffer[2093] = 21'b100000000000000000000;
 buffer[2094] = 21'b100000000000000000000;
 buffer[2095] = 21'b100000000000000000000;
 buffer[2096] = 21'b100000000000000000000;
 buffer[2097] = 21'b100000000000000000000;
 buffer[2098] = 21'b100000000000000000000;
 buffer[2099] = 21'b100000000000000000000;
 buffer[2100] = 21'b100000000000000000000;
 buffer[2101] = 21'b100000000000000000000;
 buffer[2102] = 21'b100000000000000000000;
 buffer[2103] = 21'b100000000000000000000;
 buffer[2104] = 21'b100000000000000000000;
 buffer[2105] = 21'b100000000000000000000;
 buffer[2106] = 21'b100000000000000000000;
 buffer[2107] = 21'b100000000000000000000;
 buffer[2108] = 21'b100000000000000000000;
 buffer[2109] = 21'b100000000000000000000;
 buffer[2110] = 21'b100000000000000000000;
 buffer[2111] = 21'b100000000000000000000;
 buffer[2112] = 21'b100000000000000000000;
 buffer[2113] = 21'b100000000000000000000;
 buffer[2114] = 21'b100000000000000000000;
 buffer[2115] = 21'b100000000000000000000;
 buffer[2116] = 21'b100000000000000000000;
 buffer[2117] = 21'b100000000000000000000;
 buffer[2118] = 21'b100000000000000000000;
 buffer[2119] = 21'b100000000000000000000;
 buffer[2120] = 21'b100000000000000000000;
 buffer[2121] = 21'b100000000000000000000;
 buffer[2122] = 21'b100000000000000000000;
 buffer[2123] = 21'b100000000000000000000;
 buffer[2124] = 21'b100000000000000000000;
 buffer[2125] = 21'b100000000000000000000;
 buffer[2126] = 21'b100000000000000000000;
 buffer[2127] = 21'b100000000000000000000;
 buffer[2128] = 21'b100000000000000000000;
 buffer[2129] = 21'b100000000000000000000;
 buffer[2130] = 21'b100000000000000000000;
 buffer[2131] = 21'b100000000000000000000;
 buffer[2132] = 21'b100000000000000000000;
 buffer[2133] = 21'b100000000000000000000;
 buffer[2134] = 21'b100000000000000000000;
 buffer[2135] = 21'b100000000000000000000;
 buffer[2136] = 21'b100000000000000000000;
 buffer[2137] = 21'b100000000000000000000;
 buffer[2138] = 21'b100000000000000000000;
 buffer[2139] = 21'b100000000000000000000;
 buffer[2140] = 21'b100000000000000000000;
 buffer[2141] = 21'b100000000000000000000;
 buffer[2142] = 21'b100000000000000000000;
 buffer[2143] = 21'b100000000000000000000;
 buffer[2144] = 21'b100000000000000000000;
 buffer[2145] = 21'b100000000000000000000;
 buffer[2146] = 21'b100000000000000000000;
 buffer[2147] = 21'b100000000000000000000;
 buffer[2148] = 21'b100000000000000000000;
 buffer[2149] = 21'b100000000000000000000;
 buffer[2150] = 21'b100000000000000000000;
 buffer[2151] = 21'b100000000000000000000;
 buffer[2152] = 21'b100000000000000000000;
 buffer[2153] = 21'b100000000000000000000;
 buffer[2154] = 21'b100000000000000000000;
 buffer[2155] = 21'b100000000000000000000;
 buffer[2156] = 21'b100000000000000000000;
 buffer[2157] = 21'b100000000000000000000;
 buffer[2158] = 21'b100000000000000000000;
 buffer[2159] = 21'b100000000000000000000;
 buffer[2160] = 21'b100000000000000000000;
 buffer[2161] = 21'b100000000000000000000;
 buffer[2162] = 21'b100000000000000000000;
 buffer[2163] = 21'b100000000000000000000;
 buffer[2164] = 21'b100000000000000000000;
 buffer[2165] = 21'b100000000000000000000;
 buffer[2166] = 21'b100000000000000000000;
 buffer[2167] = 21'b100000000000000000000;
 buffer[2168] = 21'b100000000000000000000;
 buffer[2169] = 21'b100000000000000000000;
 buffer[2170] = 21'b100000000000000000000;
 buffer[2171] = 21'b100000000000000000000;
 buffer[2172] = 21'b100000000000000000000;
 buffer[2173] = 21'b100000000000000000000;
 buffer[2174] = 21'b100000000000000000000;
 buffer[2175] = 21'b100000000000000000000;
 buffer[2176] = 21'b100000000000000000000;
 buffer[2177] = 21'b100000000000000000000;
 buffer[2178] = 21'b100000000000000000000;
 buffer[2179] = 21'b100000000000000000000;
 buffer[2180] = 21'b100000000000000000000;
 buffer[2181] = 21'b100000000000000000000;
 buffer[2182] = 21'b100000000000000000000;
 buffer[2183] = 21'b100000000000000000000;
 buffer[2184] = 21'b100000000000000000000;
 buffer[2185] = 21'b100000000000000000000;
 buffer[2186] = 21'b100000000000000000000;
 buffer[2187] = 21'b100000000000000000000;
 buffer[2188] = 21'b100000000000000000000;
 buffer[2189] = 21'b100000000000000000000;
 buffer[2190] = 21'b100000000000000000000;
 buffer[2191] = 21'b100000000000000000000;
 buffer[2192] = 21'b100000000000000000000;
 buffer[2193] = 21'b100000000000000000000;
 buffer[2194] = 21'b100000000000000000000;
 buffer[2195] = 21'b100000000000000000000;
 buffer[2196] = 21'b100000000000000000000;
 buffer[2197] = 21'b100000000000000000000;
 buffer[2198] = 21'b100000000000000000000;
 buffer[2199] = 21'b100000000000000000000;
 buffer[2200] = 21'b100000000000000000000;
 buffer[2201] = 21'b100000000000000000000;
 buffer[2202] = 21'b100000000000000000000;
 buffer[2203] = 21'b100000000000000000000;
 buffer[2204] = 21'b100000000000000000000;
 buffer[2205] = 21'b100000000000000000000;
 buffer[2206] = 21'b100000000000000000000;
 buffer[2207] = 21'b100000000000000000000;
 buffer[2208] = 21'b100000000000000000000;
 buffer[2209] = 21'b100000000000000000000;
 buffer[2210] = 21'b100000000000000000000;
 buffer[2211] = 21'b100000000000000000000;
 buffer[2212] = 21'b100000000000000000000;
 buffer[2213] = 21'b100000000000000000000;
 buffer[2214] = 21'b100000000000000000000;
 buffer[2215] = 21'b100000000000000000000;
 buffer[2216] = 21'b100000000000000000000;
 buffer[2217] = 21'b100000000000000000000;
 buffer[2218] = 21'b100000000000000000000;
 buffer[2219] = 21'b100000000000000000000;
 buffer[2220] = 21'b100000000000000000000;
 buffer[2221] = 21'b100000000000000000000;
 buffer[2222] = 21'b100000000000000000000;
 buffer[2223] = 21'b100000000000000000000;
 buffer[2224] = 21'b100000000000000000000;
 buffer[2225] = 21'b100000000000000000000;
 buffer[2226] = 21'b100000000000000000000;
 buffer[2227] = 21'b100000000000000000000;
 buffer[2228] = 21'b100000000000000000000;
 buffer[2229] = 21'b100000000000000000000;
 buffer[2230] = 21'b100000000000000000000;
 buffer[2231] = 21'b100000000000000000000;
 buffer[2232] = 21'b100000000000000000000;
 buffer[2233] = 21'b100000000000000000000;
 buffer[2234] = 21'b100000000000000000000;
 buffer[2235] = 21'b100000000000000000000;
 buffer[2236] = 21'b100000000000000000000;
 buffer[2237] = 21'b100000000000000000000;
 buffer[2238] = 21'b100000000000000000000;
 buffer[2239] = 21'b100000000000000000000;
 buffer[2240] = 21'b100000000000000000000;
 buffer[2241] = 21'b100000000000000000000;
 buffer[2242] = 21'b100000000000000000000;
 buffer[2243] = 21'b100000000000000000000;
 buffer[2244] = 21'b100000000000000000000;
 buffer[2245] = 21'b100000000000000000000;
 buffer[2246] = 21'b100000000000000000000;
 buffer[2247] = 21'b100000000000000000000;
 buffer[2248] = 21'b100000000000000000000;
 buffer[2249] = 21'b100000000000000000000;
 buffer[2250] = 21'b100000000000000000000;
 buffer[2251] = 21'b100000000000000000000;
 buffer[2252] = 21'b100000000000000000000;
 buffer[2253] = 21'b100000000000000000000;
 buffer[2254] = 21'b100000000000000000000;
 buffer[2255] = 21'b100000000000000000000;
 buffer[2256] = 21'b100000000000000000000;
 buffer[2257] = 21'b100000000000000000000;
 buffer[2258] = 21'b100000000000000000000;
 buffer[2259] = 21'b100000000000000000000;
 buffer[2260] = 21'b100000000000000000000;
 buffer[2261] = 21'b100000000000000000000;
 buffer[2262] = 21'b100000000000000000000;
 buffer[2263] = 21'b100000000000000000000;
 buffer[2264] = 21'b100000000000000000000;
 buffer[2265] = 21'b100000000000000000000;
 buffer[2266] = 21'b100000000000000000000;
 buffer[2267] = 21'b100000000000000000000;
 buffer[2268] = 21'b100000000000000000000;
 buffer[2269] = 21'b100000000000000000000;
 buffer[2270] = 21'b100000000000000000000;
 buffer[2271] = 21'b100000000000000000000;
 buffer[2272] = 21'b100000000000000000000;
 buffer[2273] = 21'b100000000000000000000;
 buffer[2274] = 21'b100000000000000000000;
 buffer[2275] = 21'b100000000000000000000;
 buffer[2276] = 21'b100000000000000000000;
 buffer[2277] = 21'b100000000000000000000;
 buffer[2278] = 21'b100000000000000000000;
 buffer[2279] = 21'b100000000000000000000;
 buffer[2280] = 21'b100000000000000000000;
 buffer[2281] = 21'b100000000000000000000;
 buffer[2282] = 21'b100000000000000000000;
 buffer[2283] = 21'b100000000000000000000;
 buffer[2284] = 21'b100000000000000000000;
 buffer[2285] = 21'b100000000000000000000;
 buffer[2286] = 21'b100000000000000000000;
 buffer[2287] = 21'b100000000000000000000;
 buffer[2288] = 21'b100000000000000000000;
 buffer[2289] = 21'b100000000000000000000;
 buffer[2290] = 21'b100000000000000000000;
 buffer[2291] = 21'b100000000000000000000;
 buffer[2292] = 21'b100000000000000000000;
 buffer[2293] = 21'b100000000000000000000;
 buffer[2294] = 21'b100000000000000000000;
 buffer[2295] = 21'b100000000000000000000;
 buffer[2296] = 21'b100000000000000000000;
 buffer[2297] = 21'b100000000000000000000;
 buffer[2298] = 21'b100000000000000000000;
 buffer[2299] = 21'b100000000000000000000;
 buffer[2300] = 21'b100000000000000000000;
 buffer[2301] = 21'b100000000000000000000;
 buffer[2302] = 21'b100000000000000000000;
 buffer[2303] = 21'b100000000000000000000;
 buffer[2304] = 21'b100000000000000000000;
 buffer[2305] = 21'b100000000000000000000;
 buffer[2306] = 21'b100000000000000000000;
 buffer[2307] = 21'b100000000000000000000;
 buffer[2308] = 21'b100000000000000000000;
 buffer[2309] = 21'b100000000000000000000;
 buffer[2310] = 21'b100000000000000000000;
 buffer[2311] = 21'b100000000000000000000;
 buffer[2312] = 21'b100000000000000000000;
 buffer[2313] = 21'b100000000000000000000;
 buffer[2314] = 21'b100000000000000000000;
 buffer[2315] = 21'b100000000000000000000;
 buffer[2316] = 21'b100000000000000000000;
 buffer[2317] = 21'b100000000000000000000;
 buffer[2318] = 21'b100000000000000000000;
 buffer[2319] = 21'b100000000000000000000;
 buffer[2320] = 21'b100000000000000000000;
 buffer[2321] = 21'b100000000000000000000;
 buffer[2322] = 21'b100000000000000000000;
 buffer[2323] = 21'b100000000000000000000;
 buffer[2324] = 21'b100000000000000000000;
 buffer[2325] = 21'b100000000000000000000;
 buffer[2326] = 21'b100000000000000000000;
 buffer[2327] = 21'b100000000000000000000;
 buffer[2328] = 21'b100000000000000000000;
 buffer[2329] = 21'b100000000000000000000;
 buffer[2330] = 21'b100000000000000000000;
 buffer[2331] = 21'b100000000000000000000;
 buffer[2332] = 21'b100000000000000000000;
 buffer[2333] = 21'b100000000000000000000;
 buffer[2334] = 21'b100000000000000000000;
 buffer[2335] = 21'b100000000000000000000;
 buffer[2336] = 21'b100000000000000000000;
 buffer[2337] = 21'b100000000000000000000;
 buffer[2338] = 21'b100000000000000000000;
 buffer[2339] = 21'b100000000000000000000;
 buffer[2340] = 21'b100000000000000000000;
 buffer[2341] = 21'b100000000000000000000;
 buffer[2342] = 21'b100000000000000000000;
 buffer[2343] = 21'b100000000000000000000;
 buffer[2344] = 21'b100000000000000000000;
 buffer[2345] = 21'b100000000000000000000;
 buffer[2346] = 21'b100000000000000000000;
 buffer[2347] = 21'b100000000000000000000;
 buffer[2348] = 21'b100000000000000000000;
 buffer[2349] = 21'b100000000000000000000;
 buffer[2350] = 21'b100000000000000000000;
 buffer[2351] = 21'b100000000000000000000;
 buffer[2352] = 21'b100000000000000000000;
 buffer[2353] = 21'b100000000000000000000;
 buffer[2354] = 21'b100000000000000000000;
 buffer[2355] = 21'b100000000000000000000;
 buffer[2356] = 21'b100000000000000000000;
 buffer[2357] = 21'b100000000000000000000;
 buffer[2358] = 21'b100000000000000000000;
 buffer[2359] = 21'b100000000000000000000;
 buffer[2360] = 21'b100000000000000000000;
 buffer[2361] = 21'b100000000000000000000;
 buffer[2362] = 21'b100000000000000000000;
 buffer[2363] = 21'b100000000000000000000;
 buffer[2364] = 21'b100000000000000000000;
 buffer[2365] = 21'b100000000000000000000;
 buffer[2366] = 21'b100000000000000000000;
 buffer[2367] = 21'b100000000000000000000;
 buffer[2368] = 21'b100000000000000000000;
 buffer[2369] = 21'b100000000000000000000;
 buffer[2370] = 21'b100000000000000000000;
 buffer[2371] = 21'b100000000000000000000;
 buffer[2372] = 21'b100000000000000000000;
 buffer[2373] = 21'b100000000000000000000;
 buffer[2374] = 21'b100000000000000000000;
 buffer[2375] = 21'b100000000000000000000;
 buffer[2376] = 21'b100000000000000000000;
 buffer[2377] = 21'b100000000000000000000;
 buffer[2378] = 21'b100000000000000000000;
 buffer[2379] = 21'b100000000000000000000;
 buffer[2380] = 21'b100000000000000000000;
 buffer[2381] = 21'b100000000000000000000;
 buffer[2382] = 21'b100000000000000000000;
 buffer[2383] = 21'b100000000000000000000;
 buffer[2384] = 21'b100000000000000000000;
 buffer[2385] = 21'b100000000000000000000;
 buffer[2386] = 21'b100000000000000000000;
 buffer[2387] = 21'b100000000000000000000;
 buffer[2388] = 21'b100000000000000000000;
 buffer[2389] = 21'b100000000000000000000;
 buffer[2390] = 21'b100000000000000000000;
 buffer[2391] = 21'b100000000000000000000;
 buffer[2392] = 21'b100000000000000000000;
 buffer[2393] = 21'b100000000000000000000;
 buffer[2394] = 21'b100000000000000000000;
 buffer[2395] = 21'b100000000000000000000;
 buffer[2396] = 21'b100000000000000000000;
 buffer[2397] = 21'b100000000000000000000;
 buffer[2398] = 21'b100000000000000000000;
 buffer[2399] = 21'b100000000000000000000;
end

endmodule

module M_character_map (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_tpu_x,
in_tpu_y,
in_tpu_character,
in_tpu_foreground,
in_tpu_background,
in_tpu_write,
out_pix_red,
out_pix_green,
out_pix_blue,
out_character_map_display,
out_tpu_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [6:0] in_tpu_x;
input  [4:0] in_tpu_y;
input  [7:0] in_tpu_character;
input  [5:0] in_tpu_foreground;
input  [6:0] in_tpu_background;
input  [2:0] in_tpu_write;
output  [1:0] out_pix_red;
output  [1:0] out_pix_green;
output  [1:0] out_pix_blue;
output  [0:0] out_character_map_display;
output  [0:0] out_tpu_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [7:0] _w_mem_characterGenerator8x16_rdata;
wire  [20:0] _w_mem_charactermap_rdata0;
wire  [7:0] _w_xcharacterpos;
wire  [11:0] _w_ycharacterpos;
wire  [2:0] _w_xincharacter;
wire  [3:0] _w_yincharacter;
wire  [0:0] _w_characterpixel;

reg  [11:0] _d_characterGenerator8x16_addr;
reg  [11:0] _q_characterGenerator8x16_addr;
reg  [11:0] _d_charactermap_addr0;
reg  [11:0] _q_charactermap_addr0;
reg  [0:0] _d_charactermap_wenable1;
reg  [0:0] _q_charactermap_wenable1;
reg  [20:0] _d_charactermap_wdata1;
reg  [20:0] _q_charactermap_wdata1;
reg  [11:0] _d_charactermap_addr1;
reg  [11:0] _q_charactermap_addr1;
reg  [6:0] _d_tpu_active_x;
reg  [6:0] _q_tpu_active_x;
reg  [4:0] _d_tpu_active_y;
reg  [4:0] _q_tpu_active_y;
reg  [11:0] _d_tpu_cs_addr;
reg  [11:0] _q_tpu_cs_addr;
reg  [1:0] _d_pix_red,_q_pix_red;
reg  [1:0] _d_pix_green,_q_pix_green;
reg  [1:0] _d_pix_blue,_q_pix_blue;
reg  [0:0] _d_character_map_display,_q_character_map_display;
reg  [0:0] _d_tpu_active,_q_tpu_active;
reg  [2:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_character_map_display = _d_character_map_display;
assign out_tpu_active = _q_tpu_active;
assign out_done = (_q_index == 5);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_characterGenerator8x16_addr <= 0;
_q_charactermap_addr0 <= 0;
_q_charactermap_wenable1 <= 0;
_q_charactermap_wdata1 <= 0;
_q_charactermap_addr1 <= 0;
_q_tpu_active_x <= 0;
_q_tpu_active_y <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_characterGenerator8x16_addr <= _d_characterGenerator8x16_addr;
_q_charactermap_addr0 <= _d_charactermap_addr0;
_q_charactermap_wenable1 <= _d_charactermap_wenable1;
_q_charactermap_wdata1 <= _d_charactermap_wdata1;
_q_charactermap_addr1 <= _d_charactermap_addr1;
_q_tpu_active_x <= _d_tpu_active_x;
_q_tpu_active_y <= _d_tpu_active_y;
_q_tpu_cs_addr <= _d_tpu_cs_addr;
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_character_map_display <= _d_character_map_display;
_q_tpu_active <= _d_tpu_active;
_q_index <= _d_index;
  end
end


M_character_map_mem_characterGenerator8x16 __mem__characterGenerator8x16(
.clock(clock),
.in_characterGenerator8x16_addr(_d_characterGenerator8x16_addr),
.out_characterGenerator8x16_rdata(_w_mem_characterGenerator8x16_rdata)
);
M_character_map_mem_charactermap __mem__charactermap(
.clock0(clock),
.clock1(clock),
.in_charactermap_addr0(_d_charactermap_addr0),
.in_charactermap_wenable1(_d_charactermap_wenable1),
.in_charactermap_wdata1(_d_charactermap_wdata1),
.in_charactermap_addr1(_d_charactermap_addr1),
.out_charactermap_rdata0(_w_mem_charactermap_rdata0)
);

assign _w_characterpixel = _w_mem_characterGenerator8x16_rdata[7-_w_xincharacter+:1];
assign _w_yincharacter = (in_pix_y)&15;
assign _w_ycharacterpos = ((in_pix_vblank?0:in_pix_y)>>4)*80;
assign _w_xincharacter = (in_pix_x)&7;
assign _w_xcharacterpos = (in_pix_active?in_pix_x+2:0)>>3;

always @* begin
_d_characterGenerator8x16_addr = _q_characterGenerator8x16_addr;
_d_charactermap_addr0 = _q_charactermap_addr0;
_d_charactermap_wenable1 = _q_charactermap_wenable1;
_d_charactermap_wdata1 = _q_charactermap_wdata1;
_d_charactermap_addr1 = _q_charactermap_addr1;
_d_tpu_active_x = _q_tpu_active_x;
_d_tpu_active_y = _q_tpu_active_y;
_d_tpu_cs_addr = _q_tpu_cs_addr;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_character_map_display = _q_character_map_display;
_d_tpu_active = _q_tpu_active;
_d_index = _q_index;
// _always_pre
_d_charactermap_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_charactermap_wenable1 = 1;
_d_characterGenerator8x16_addr = _w_mem_charactermap_rdata0[0+:8]*16+_w_yincharacter;
_d_character_map_display = in_pix_active&&((_w_characterpixel)||(~_w_mem_charactermap_rdata0[20+:1]));
_d_pix_red = _w_characterpixel?_w_mem_charactermap_rdata0[12+:2]:_w_mem_charactermap_rdata0[18+:2];
_d_pix_green = _w_characterpixel?_w_mem_charactermap_rdata0[10+:2]:_w_mem_charactermap_rdata0[16+:2];
_d_pix_blue = _w_characterpixel?_w_mem_charactermap_rdata0[8+:2]:_w_mem_charactermap_rdata0[14+:2];
_d_index = 5;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_characterGenerator8x16_addr = 0;
_d_charactermap_addr0 = 0;
_d_charactermap_wenable1 = 0;
_d_charactermap_wdata1 = 0;
_d_charactermap_addr1 = 0;
_d_tpu_active_x = 0;
_d_tpu_active_y = 0;
// --
_d_charactermap_addr1 = 0;
_d_charactermap_wdata1 = {1'b1,6'b0,6'b0,8'b0};
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (_q_tpu_active)
  0: begin
// __block_6_case
// __block_7
  case (in_tpu_write)
  1: begin
// __block_9_case
// __block_10
_d_tpu_active_x = in_tpu_x;
_d_tpu_active_y = in_tpu_y;
// __block_11
  end
  2: begin
// __block_12_case
// __block_13
_d_charactermap_addr1 = _q_tpu_active_x+_q_tpu_active_y*80;
_d_charactermap_wdata1 = {in_tpu_background,in_tpu_foreground,in_tpu_character};
_d_tpu_active_y = (_q_tpu_active_x==79)?(_q_tpu_active_y==29)?0:_q_tpu_active_y+1:_q_tpu_active_y;
_d_tpu_active_x = (_q_tpu_active_x==79)?0:_q_tpu_active_x+1;
// __block_14
  end
  3: begin
// __block_15_case
// __block_16
_d_tpu_active_x = 0;
_d_tpu_active_y = 0;
_d_tpu_active = 1;
_d_tpu_cs_addr = 0;
_d_charactermap_wdata1 = {1'b1,6'b0,6'b0,8'b0};
// __block_17
  end
endcase
// __block_8
// __block_18
_d_index = 1;
  end
  1: begin
// __block_19_case
// __block_20
_d_index = 3;
  end
endcase
end else begin
_d_index = 2;
end
end
3: begin
// __while__block_21
if (_q_tpu_cs_addr<2400) begin
// __block_22
// __block_24
_d_charactermap_addr1 = _q_tpu_cs_addr;
_d_tpu_cs_addr = _q_tpu_cs_addr+1;
// __block_25
_d_index = 3;
end else begin
_d_index = 4;
end
end
2: begin
// __block_3
_d_index = 5;
end
4: begin
// __block_26
_d_tpu_active = 0;
// __block_27
_d_index = 1;
end
5: begin // end of character_map
end
default: begin 
_d_index = 5;
 end
endcase
end
endmodule


module M_bitmap #(
parameter BITMAP_ADDR0_WIDTH=1,parameter BITMAP_ADDR0_SIGNED=0,parameter BITMAP_ADDR0_INIT=0,
parameter BITMAP_RDATA0_WIDTH=1,parameter BITMAP_RDATA0_SIGNED=0,parameter BITMAP_RDATA0_INIT=0
) (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_bitmap_write_offset,
in_bitmap_x_read,
in_bitmap_y_read,
in_bitmap_rdata0,
out_pix_red,
out_pix_green,
out_pix_blue,
out_bitmap_display,
out_x_offset,
out_y_offset,
out_bitmap_colour_read,
out_bitmap_addr0,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [2:0] in_bitmap_write_offset;
input signed [15:0] in_bitmap_x_read;
input signed [15:0] in_bitmap_y_read;
input  [BITMAP_RDATA0_WIDTH-1:0] in_bitmap_rdata0;
output  [1:0] out_pix_red;
output  [1:0] out_pix_green;
output  [1:0] out_pix_blue;
output  [0:0] out_bitmap_display;
output  [9:0] out_x_offset;
output  [9:0] out_y_offset;
output  [6:0] out_bitmap_colour_read;
output  [BITMAP_ADDR0_WIDTH-1:0] out_bitmap_addr0;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [9:0] _w_x_plus_one;
wire  [9:0] _w_y_line;
wire  [9:0] _w_x_pixel;

reg  [1:0] _d_pix_red,_q_pix_red;
reg  [1:0] _d_pix_green,_q_pix_green;
reg  [1:0] _d_pix_blue,_q_pix_blue;
reg  [0:0] _d_bitmap_display,_q_bitmap_display;
reg  [9:0] _d_x_offset,_q_x_offset;
reg  [9:0] _d_y_offset,_q_y_offset;
reg  [6:0] _d_bitmap_colour_read,_q_bitmap_colour_read;
reg  [BITMAP_ADDR0_WIDTH-1:0] _d_bitmap_addr0,_q_bitmap_addr0;
reg  [1:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_bitmap_display = _d_bitmap_display;
assign out_x_offset = _q_x_offset;
assign out_y_offset = _q_y_offset;
assign out_bitmap_colour_read = _q_bitmap_colour_read;
assign out_bitmap_addr0 = _d_bitmap_addr0;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_bitmap_addr0 <= BITMAP_ADDR0_INIT;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_bitmap_display <= _d_bitmap_display;
_q_x_offset <= _d_x_offset;
_q_y_offset <= _d_y_offset;
_q_bitmap_colour_read <= _d_bitmap_colour_read;
_q_bitmap_addr0 <= _d_bitmap_addr0;
_q_index <= _d_index;
  end
end



assign _w_x_pixel = in_pix_active?_w_x_plus_one:_d_x_offset;
assign _w_y_line = in_pix_vblank?_d_y_offset:((in_pix_y+_d_y_offset)>479?(in_pix_y+_d_y_offset)-479:(in_pix_y+_d_y_offset));
assign _w_x_plus_one = (in_pix_x+_d_x_offset+1)>639?(in_pix_x+_d_x_offset+1)-639:(in_pix_x+_d_x_offset+1);

always @* begin
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_bitmap_display = _q_bitmap_display;
_d_x_offset = _q_x_offset;
_d_y_offset = _q_y_offset;
_d_bitmap_colour_read = _q_bitmap_colour_read;
_d_bitmap_addr0 = _q_bitmap_addr0;
_d_index = _q_index;
// _always_pre
_d_bitmap_colour_read = (in_pix_x==in_bitmap_x_read)&&(in_pix_y==in_bitmap_y_read)?in_bitmap_rdata0:_q_bitmap_colour_read;
_d_bitmap_addr0 = _w_x_pixel+(_w_y_line*640);
_d_bitmap_display = in_pix_active&&~in_bitmap_rdata0[6+:1];
_d_pix_red = in_bitmap_rdata0[4+:2];
_d_pix_green = in_bitmap_rdata0[2+:2];
_d_pix_blue = in_bitmap_rdata0[0+:2];
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (in_bitmap_write_offset)
  1: begin
// __block_6_case
// __block_7
_d_x_offset = (_q_x_offset==639)?0:_q_x_offset+1;
// __block_8
  end
  2: begin
// __block_9_case
// __block_10
_d_y_offset = (_q_y_offset==479)?0:_q_y_offset+1;
// __block_11
  end
  3: begin
// __block_12_case
// __block_13
_d_x_offset = (_q_x_offset==0)?639:_q_x_offset-1;
// __block_14
  end
  4: begin
// __block_15_case
// __block_16
_d_y_offset = (_q_y_offset==0)?479:_q_y_offset-1;
// __block_17
  end
  5: begin
// __block_18_case
// __block_19
_d_x_offset = 0;
_d_y_offset = 0;
// __block_20
  end
endcase
// __block_5
// __block_21
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of bitmap
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_bitmapwriter #(
parameter BITMAP_ADDR1_WIDTH=1,parameter BITMAP_ADDR1_SIGNED=0,parameter BITMAP_ADDR1_INIT=0,
parameter BITMAP_WENABLE1_WIDTH=1,parameter BITMAP_WENABLE1_SIGNED=0,parameter BITMAP_WENABLE1_INIT=0,
parameter BITMAP_WDATA1_WIDTH=1,parameter BITMAP_WDATA1_SIGNED=0,parameter BITMAP_WDATA1_INIT=0
) (
in_bitmap_x_write,
in_bitmap_y_write,
in_bitmap_colour_write,
in_bitmap_write,
in_x_offset,
in_y_offset,
out_bitmap_addr1,
out_bitmap_wenable1,
out_bitmap_wdata1,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_bitmap_x_write;
input signed [10:0] in_bitmap_y_write;
input  [6:0] in_bitmap_colour_write;
input  [0:0] in_bitmap_write;
input  [9:0] in_x_offset;
input  [9:0] in_y_offset;
output  [BITMAP_ADDR1_WIDTH-1:0] out_bitmap_addr1;
output  [BITMAP_WENABLE1_WIDTH-1:0] out_bitmap_wenable1;
output  [BITMAP_WDATA1_WIDTH-1:0] out_bitmap_wdata1;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [9:0] _w_x_write_pixel;
wire  [9:0] _w_y_write_pixel;
wire  [0:0] _w_write_pixel;

reg  [BITMAP_ADDR1_WIDTH-1:0] _d_bitmap_addr1,_q_bitmap_addr1;
reg  [BITMAP_WENABLE1_WIDTH-1:0] _d_bitmap_wenable1,_q_bitmap_wenable1;
reg  [BITMAP_WDATA1_WIDTH-1:0] _d_bitmap_wdata1,_q_bitmap_wdata1;
reg  [1:0] _d_index,_q_index;
assign out_bitmap_addr1 = _d_bitmap_addr1;
assign out_bitmap_wenable1 = _d_bitmap_wenable1;
assign out_bitmap_wdata1 = _d_bitmap_wdata1;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_bitmap_addr1 <= BITMAP_ADDR1_INIT;
_q_bitmap_wenable1 <= BITMAP_WENABLE1_INIT;
_q_bitmap_wdata1 <= BITMAP_WDATA1_INIT;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_bitmap_addr1 <= _d_bitmap_addr1;
_q_bitmap_wenable1 <= _d_bitmap_wenable1;
_q_bitmap_wdata1 <= _d_bitmap_wdata1;
_q_index <= _d_index;
  end
end



assign _w_write_pixel = (in_bitmap_x_write>=0)&&(in_bitmap_x_write<640)&&(in_bitmap_y_write>=0)&&(in_bitmap_y_write<=479)&&in_bitmap_write;
assign _w_y_write_pixel = (in_bitmap_y_write+in_y_offset)>479?(in_bitmap_y_write+in_y_offset)-479:(in_bitmap_y_write+in_y_offset);
assign _w_x_write_pixel = (in_bitmap_x_write+in_x_offset)>639?(in_bitmap_x_write+in_x_offset)-639:(in_bitmap_x_write+in_x_offset);

always @* begin
_d_bitmap_addr1 = _q_bitmap_addr1;
_d_bitmap_wenable1 = _q_bitmap_wenable1;
_d_bitmap_wdata1 = _q_bitmap_wdata1;
_d_index = _q_index;
// _always_pre
_d_bitmap_wenable1 = 1;
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (_w_write_pixel==1) begin
// __block_5
// __block_7
_d_bitmap_addr1 = _w_x_write_pixel+_w_y_write_pixel*640;
_d_bitmap_wdata1 = in_bitmap_colour_write;
// __block_8
end else begin
// __block_6
end
// __block_9
// __block_10
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of bitmapwriter
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_gpu_mem_blit1tilemap(
input      [8:0]                in_blit1tilemap_addr0,
output reg  [15:0]     out_blit1tilemap_rdata0,
output reg  [15:0]     out_blit1tilemap_rdata1,
input      [0:0]             in_blit1tilemap_wenable1,
input      [15:0]                 in_blit1tilemap_wdata1,
input      [8:0]                in_blit1tilemap_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[511:0];
always @(posedge clock0) begin
  out_blit1tilemap_rdata0 <= buffer[in_blit1tilemap_addr0];
end
always @(posedge clock1) begin
  if (in_blit1tilemap_wenable1) begin
    buffer[in_blit1tilemap_addr1] <= in_blit1tilemap_wdata1;
  end
end

endmodule

module M_gpu_mem_characterGenerator8x8(
input      [10:0]                in_characterGenerator8x8_addr0,
output reg  [7:0]     out_characterGenerator8x8_rdata0,
output reg  [7:0]     out_characterGenerator8x8_rdata1,
input      [0:0]             in_characterGenerator8x8_wenable1,
input      [7:0]                 in_characterGenerator8x8_wdata1,
input      [10:0]                in_characterGenerator8x8_addr1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2047:0];
always @(posedge clock0) begin
  out_characterGenerator8x8_rdata0 <= buffer[in_characterGenerator8x8_addr0];
end
always @(posedge clock1) begin
  if (in_characterGenerator8x8_wenable1) begin
    buffer[in_characterGenerator8x8_addr1] <= in_characterGenerator8x8_wdata1;
  end
end
initial begin
 buffer[0] = 8'h00;
 buffer[1] = 8'h00;
 buffer[2] = 8'h00;
 buffer[3] = 8'h00;
 buffer[4] = 8'h00;
 buffer[5] = 8'h00;
 buffer[6] = 8'h00;
 buffer[7] = 8'h00;
 buffer[8] = 8'h7e;
 buffer[9] = 8'h81;
 buffer[10] = 8'ha5;
 buffer[11] = 8'h81;
 buffer[12] = 8'hbd;
 buffer[13] = 8'h99;
 buffer[14] = 8'h81;
 buffer[15] = 8'h7e;
 buffer[16] = 8'h7e;
 buffer[17] = 8'hff;
 buffer[18] = 8'hdb;
 buffer[19] = 8'hff;
 buffer[20] = 8'hc3;
 buffer[21] = 8'he7;
 buffer[22] = 8'hff;
 buffer[23] = 8'h7e;
 buffer[24] = 8'h6c;
 buffer[25] = 8'hfe;
 buffer[26] = 8'hfe;
 buffer[27] = 8'hfe;
 buffer[28] = 8'h7c;
 buffer[29] = 8'h38;
 buffer[30] = 8'h10;
 buffer[31] = 8'h00;
 buffer[32] = 8'h10;
 buffer[33] = 8'h38;
 buffer[34] = 8'h7c;
 buffer[35] = 8'hfe;
 buffer[36] = 8'h7c;
 buffer[37] = 8'h38;
 buffer[38] = 8'h10;
 buffer[39] = 8'h00;
 buffer[40] = 8'h38;
 buffer[41] = 8'h7c;
 buffer[42] = 8'h38;
 buffer[43] = 8'hfe;
 buffer[44] = 8'hfe;
 buffer[45] = 8'h7c;
 buffer[46] = 8'h38;
 buffer[47] = 8'h7c;
 buffer[48] = 8'h10;
 buffer[49] = 8'h10;
 buffer[50] = 8'h38;
 buffer[51] = 8'h7c;
 buffer[52] = 8'hfe;
 buffer[53] = 8'h7c;
 buffer[54] = 8'h38;
 buffer[55] = 8'h7c;
 buffer[56] = 8'h00;
 buffer[57] = 8'h00;
 buffer[58] = 8'h18;
 buffer[59] = 8'h3c;
 buffer[60] = 8'h3c;
 buffer[61] = 8'h18;
 buffer[62] = 8'h00;
 buffer[63] = 8'h00;
 buffer[64] = 8'hff;
 buffer[65] = 8'hff;
 buffer[66] = 8'he7;
 buffer[67] = 8'hc3;
 buffer[68] = 8'hc3;
 buffer[69] = 8'he7;
 buffer[70] = 8'hff;
 buffer[71] = 8'hff;
 buffer[72] = 8'h00;
 buffer[73] = 8'h3c;
 buffer[74] = 8'h66;
 buffer[75] = 8'h42;
 buffer[76] = 8'h42;
 buffer[77] = 8'h66;
 buffer[78] = 8'h3c;
 buffer[79] = 8'h00;
 buffer[80] = 8'hff;
 buffer[81] = 8'hc3;
 buffer[82] = 8'h99;
 buffer[83] = 8'hbd;
 buffer[84] = 8'hbd;
 buffer[85] = 8'h99;
 buffer[86] = 8'hc3;
 buffer[87] = 8'hff;
 buffer[88] = 8'h0f;
 buffer[89] = 8'h07;
 buffer[90] = 8'h0f;
 buffer[91] = 8'h7d;
 buffer[92] = 8'hcc;
 buffer[93] = 8'hcc;
 buffer[94] = 8'hcc;
 buffer[95] = 8'h78;
 buffer[96] = 8'h3c;
 buffer[97] = 8'h66;
 buffer[98] = 8'h66;
 buffer[99] = 8'h66;
 buffer[100] = 8'h3c;
 buffer[101] = 8'h18;
 buffer[102] = 8'h7e;
 buffer[103] = 8'h18;
 buffer[104] = 8'h3f;
 buffer[105] = 8'h33;
 buffer[106] = 8'h3f;
 buffer[107] = 8'h30;
 buffer[108] = 8'h30;
 buffer[109] = 8'h70;
 buffer[110] = 8'hf0;
 buffer[111] = 8'he0;
 buffer[112] = 8'h7f;
 buffer[113] = 8'h63;
 buffer[114] = 8'h7f;
 buffer[115] = 8'h63;
 buffer[116] = 8'h63;
 buffer[117] = 8'h67;
 buffer[118] = 8'he6;
 buffer[119] = 8'hc0;
 buffer[120] = 8'h99;
 buffer[121] = 8'h5a;
 buffer[122] = 8'h3c;
 buffer[123] = 8'he7;
 buffer[124] = 8'he7;
 buffer[125] = 8'h3c;
 buffer[126] = 8'h5a;
 buffer[127] = 8'h99;
 buffer[128] = 8'h80;
 buffer[129] = 8'he0;
 buffer[130] = 8'hf8;
 buffer[131] = 8'hfe;
 buffer[132] = 8'hf8;
 buffer[133] = 8'he0;
 buffer[134] = 8'h80;
 buffer[135] = 8'h00;
 buffer[136] = 8'h02;
 buffer[137] = 8'h0e;
 buffer[138] = 8'h3e;
 buffer[139] = 8'hfe;
 buffer[140] = 8'h3e;
 buffer[141] = 8'h0e;
 buffer[142] = 8'h02;
 buffer[143] = 8'h00;
 buffer[144] = 8'h18;
 buffer[145] = 8'h3c;
 buffer[146] = 8'h7e;
 buffer[147] = 8'h18;
 buffer[148] = 8'h18;
 buffer[149] = 8'h7e;
 buffer[150] = 8'h3c;
 buffer[151] = 8'h18;
 buffer[152] = 8'h66;
 buffer[153] = 8'h66;
 buffer[154] = 8'h66;
 buffer[155] = 8'h66;
 buffer[156] = 8'h66;
 buffer[157] = 8'h00;
 buffer[158] = 8'h66;
 buffer[159] = 8'h00;
 buffer[160] = 8'h7f;
 buffer[161] = 8'hdb;
 buffer[162] = 8'hdb;
 buffer[163] = 8'h7b;
 buffer[164] = 8'h1b;
 buffer[165] = 8'h1b;
 buffer[166] = 8'h1b;
 buffer[167] = 8'h00;
 buffer[168] = 8'h3e;
 buffer[169] = 8'h63;
 buffer[170] = 8'h38;
 buffer[171] = 8'h6c;
 buffer[172] = 8'h6c;
 buffer[173] = 8'h38;
 buffer[174] = 8'hcc;
 buffer[175] = 8'h78;
 buffer[176] = 8'h00;
 buffer[177] = 8'h00;
 buffer[178] = 8'h00;
 buffer[179] = 8'h00;
 buffer[180] = 8'h7e;
 buffer[181] = 8'h7e;
 buffer[182] = 8'h7e;
 buffer[183] = 8'h00;
 buffer[184] = 8'h18;
 buffer[185] = 8'h3c;
 buffer[186] = 8'h7e;
 buffer[187] = 8'h18;
 buffer[188] = 8'h7e;
 buffer[189] = 8'h3c;
 buffer[190] = 8'h18;
 buffer[191] = 8'hff;
 buffer[192] = 8'h18;
 buffer[193] = 8'h3c;
 buffer[194] = 8'h7e;
 buffer[195] = 8'h18;
 buffer[196] = 8'h18;
 buffer[197] = 8'h18;
 buffer[198] = 8'h18;
 buffer[199] = 8'h00;
 buffer[200] = 8'h18;
 buffer[201] = 8'h18;
 buffer[202] = 8'h18;
 buffer[203] = 8'h18;
 buffer[204] = 8'h7e;
 buffer[205] = 8'h3c;
 buffer[206] = 8'h18;
 buffer[207] = 8'h00;
 buffer[208] = 8'h00;
 buffer[209] = 8'h18;
 buffer[210] = 8'h0c;
 buffer[211] = 8'hfe;
 buffer[212] = 8'h0c;
 buffer[213] = 8'h18;
 buffer[214] = 8'h00;
 buffer[215] = 8'h00;
 buffer[216] = 8'h00;
 buffer[217] = 8'h30;
 buffer[218] = 8'h60;
 buffer[219] = 8'hfe;
 buffer[220] = 8'h60;
 buffer[221] = 8'h30;
 buffer[222] = 8'h00;
 buffer[223] = 8'h00;
 buffer[224] = 8'h00;
 buffer[225] = 8'h00;
 buffer[226] = 8'hc0;
 buffer[227] = 8'hc0;
 buffer[228] = 8'hc0;
 buffer[229] = 8'hfe;
 buffer[230] = 8'h00;
 buffer[231] = 8'h00;
 buffer[232] = 8'h00;
 buffer[233] = 8'h24;
 buffer[234] = 8'h66;
 buffer[235] = 8'hff;
 buffer[236] = 8'h66;
 buffer[237] = 8'h24;
 buffer[238] = 8'h00;
 buffer[239] = 8'h00;
 buffer[240] = 8'h00;
 buffer[241] = 8'h18;
 buffer[242] = 8'h3c;
 buffer[243] = 8'h7e;
 buffer[244] = 8'hff;
 buffer[245] = 8'hff;
 buffer[246] = 8'h00;
 buffer[247] = 8'h00;
 buffer[248] = 8'h00;
 buffer[249] = 8'hff;
 buffer[250] = 8'hff;
 buffer[251] = 8'h7e;
 buffer[252] = 8'h3c;
 buffer[253] = 8'h18;
 buffer[254] = 8'h00;
 buffer[255] = 8'h00;
 buffer[256] = 8'h00;
 buffer[257] = 8'h00;
 buffer[258] = 8'h00;
 buffer[259] = 8'h00;
 buffer[260] = 8'h00;
 buffer[261] = 8'h00;
 buffer[262] = 8'h00;
 buffer[263] = 8'h00;
 buffer[264] = 8'h30;
 buffer[265] = 8'h78;
 buffer[266] = 8'h78;
 buffer[267] = 8'h30;
 buffer[268] = 8'h30;
 buffer[269] = 8'h00;
 buffer[270] = 8'h30;
 buffer[271] = 8'h00;
 buffer[272] = 8'h6c;
 buffer[273] = 8'h6c;
 buffer[274] = 8'h6c;
 buffer[275] = 8'h00;
 buffer[276] = 8'h00;
 buffer[277] = 8'h00;
 buffer[278] = 8'h00;
 buffer[279] = 8'h00;
 buffer[280] = 8'h6c;
 buffer[281] = 8'h6c;
 buffer[282] = 8'hfe;
 buffer[283] = 8'h6c;
 buffer[284] = 8'hfe;
 buffer[285] = 8'h6c;
 buffer[286] = 8'h6c;
 buffer[287] = 8'h00;
 buffer[288] = 8'h30;
 buffer[289] = 8'h7c;
 buffer[290] = 8'hc0;
 buffer[291] = 8'h78;
 buffer[292] = 8'h0c;
 buffer[293] = 8'hf8;
 buffer[294] = 8'h30;
 buffer[295] = 8'h00;
 buffer[296] = 8'h00;
 buffer[297] = 8'hc6;
 buffer[298] = 8'hcc;
 buffer[299] = 8'h18;
 buffer[300] = 8'h30;
 buffer[301] = 8'h66;
 buffer[302] = 8'hc6;
 buffer[303] = 8'h00;
 buffer[304] = 8'h38;
 buffer[305] = 8'h6c;
 buffer[306] = 8'h38;
 buffer[307] = 8'h76;
 buffer[308] = 8'hdc;
 buffer[309] = 8'hcc;
 buffer[310] = 8'h76;
 buffer[311] = 8'h00;
 buffer[312] = 8'h60;
 buffer[313] = 8'h60;
 buffer[314] = 8'hc0;
 buffer[315] = 8'h00;
 buffer[316] = 8'h00;
 buffer[317] = 8'h00;
 buffer[318] = 8'h00;
 buffer[319] = 8'h00;
 buffer[320] = 8'h18;
 buffer[321] = 8'h30;
 buffer[322] = 8'h60;
 buffer[323] = 8'h60;
 buffer[324] = 8'h60;
 buffer[325] = 8'h30;
 buffer[326] = 8'h18;
 buffer[327] = 8'h00;
 buffer[328] = 8'h60;
 buffer[329] = 8'h30;
 buffer[330] = 8'h18;
 buffer[331] = 8'h18;
 buffer[332] = 8'h18;
 buffer[333] = 8'h30;
 buffer[334] = 8'h60;
 buffer[335] = 8'h00;
 buffer[336] = 8'h00;
 buffer[337] = 8'h66;
 buffer[338] = 8'h3c;
 buffer[339] = 8'hff;
 buffer[340] = 8'h3c;
 buffer[341] = 8'h66;
 buffer[342] = 8'h00;
 buffer[343] = 8'h00;
 buffer[344] = 8'h00;
 buffer[345] = 8'h30;
 buffer[346] = 8'h30;
 buffer[347] = 8'hfc;
 buffer[348] = 8'h30;
 buffer[349] = 8'h30;
 buffer[350] = 8'h00;
 buffer[351] = 8'h00;
 buffer[352] = 8'h00;
 buffer[353] = 8'h00;
 buffer[354] = 8'h00;
 buffer[355] = 8'h00;
 buffer[356] = 8'h00;
 buffer[357] = 8'h30;
 buffer[358] = 8'h30;
 buffer[359] = 8'h60;
 buffer[360] = 8'h00;
 buffer[361] = 8'h00;
 buffer[362] = 8'h00;
 buffer[363] = 8'hfc;
 buffer[364] = 8'h00;
 buffer[365] = 8'h00;
 buffer[366] = 8'h00;
 buffer[367] = 8'h00;
 buffer[368] = 8'h00;
 buffer[369] = 8'h00;
 buffer[370] = 8'h00;
 buffer[371] = 8'h00;
 buffer[372] = 8'h00;
 buffer[373] = 8'h30;
 buffer[374] = 8'h30;
 buffer[375] = 8'h00;
 buffer[376] = 8'h06;
 buffer[377] = 8'h0c;
 buffer[378] = 8'h18;
 buffer[379] = 8'h30;
 buffer[380] = 8'h60;
 buffer[381] = 8'hc0;
 buffer[382] = 8'h80;
 buffer[383] = 8'h00;
 buffer[384] = 8'h7c;
 buffer[385] = 8'hc6;
 buffer[386] = 8'hce;
 buffer[387] = 8'hde;
 buffer[388] = 8'hf6;
 buffer[389] = 8'he6;
 buffer[390] = 8'h7c;
 buffer[391] = 8'h00;
 buffer[392] = 8'h30;
 buffer[393] = 8'h70;
 buffer[394] = 8'h30;
 buffer[395] = 8'h30;
 buffer[396] = 8'h30;
 buffer[397] = 8'h30;
 buffer[398] = 8'hfc;
 buffer[399] = 8'h00;
 buffer[400] = 8'h78;
 buffer[401] = 8'hcc;
 buffer[402] = 8'h0c;
 buffer[403] = 8'h38;
 buffer[404] = 8'h60;
 buffer[405] = 8'hcc;
 buffer[406] = 8'hfc;
 buffer[407] = 8'h00;
 buffer[408] = 8'h78;
 buffer[409] = 8'hcc;
 buffer[410] = 8'h0c;
 buffer[411] = 8'h38;
 buffer[412] = 8'h0c;
 buffer[413] = 8'hcc;
 buffer[414] = 8'h78;
 buffer[415] = 8'h00;
 buffer[416] = 8'h1c;
 buffer[417] = 8'h3c;
 buffer[418] = 8'h6c;
 buffer[419] = 8'hcc;
 buffer[420] = 8'hfe;
 buffer[421] = 8'h0c;
 buffer[422] = 8'h1e;
 buffer[423] = 8'h00;
 buffer[424] = 8'hfc;
 buffer[425] = 8'hc0;
 buffer[426] = 8'hf8;
 buffer[427] = 8'h0c;
 buffer[428] = 8'h0c;
 buffer[429] = 8'hcc;
 buffer[430] = 8'h78;
 buffer[431] = 8'h00;
 buffer[432] = 8'h38;
 buffer[433] = 8'h60;
 buffer[434] = 8'hc0;
 buffer[435] = 8'hf8;
 buffer[436] = 8'hcc;
 buffer[437] = 8'hcc;
 buffer[438] = 8'h78;
 buffer[439] = 8'h00;
 buffer[440] = 8'hfc;
 buffer[441] = 8'hcc;
 buffer[442] = 8'h0c;
 buffer[443] = 8'h18;
 buffer[444] = 8'h30;
 buffer[445] = 8'h30;
 buffer[446] = 8'h30;
 buffer[447] = 8'h00;
 buffer[448] = 8'h78;
 buffer[449] = 8'hcc;
 buffer[450] = 8'hcc;
 buffer[451] = 8'h78;
 buffer[452] = 8'hcc;
 buffer[453] = 8'hcc;
 buffer[454] = 8'h78;
 buffer[455] = 8'h00;
 buffer[456] = 8'h78;
 buffer[457] = 8'hcc;
 buffer[458] = 8'hcc;
 buffer[459] = 8'h7c;
 buffer[460] = 8'h0c;
 buffer[461] = 8'h18;
 buffer[462] = 8'h70;
 buffer[463] = 8'h00;
 buffer[464] = 8'h00;
 buffer[465] = 8'h30;
 buffer[466] = 8'h30;
 buffer[467] = 8'h00;
 buffer[468] = 8'h00;
 buffer[469] = 8'h30;
 buffer[470] = 8'h30;
 buffer[471] = 8'h00;
 buffer[472] = 8'h00;
 buffer[473] = 8'h30;
 buffer[474] = 8'h30;
 buffer[475] = 8'h00;
 buffer[476] = 8'h00;
 buffer[477] = 8'h30;
 buffer[478] = 8'h30;
 buffer[479] = 8'h60;
 buffer[480] = 8'h18;
 buffer[481] = 8'h30;
 buffer[482] = 8'h60;
 buffer[483] = 8'hc0;
 buffer[484] = 8'h60;
 buffer[485] = 8'h30;
 buffer[486] = 8'h18;
 buffer[487] = 8'h00;
 buffer[488] = 8'h00;
 buffer[489] = 8'h00;
 buffer[490] = 8'hfc;
 buffer[491] = 8'h00;
 buffer[492] = 8'h00;
 buffer[493] = 8'hfc;
 buffer[494] = 8'h00;
 buffer[495] = 8'h00;
 buffer[496] = 8'h60;
 buffer[497] = 8'h30;
 buffer[498] = 8'h18;
 buffer[499] = 8'h0c;
 buffer[500] = 8'h18;
 buffer[501] = 8'h30;
 buffer[502] = 8'h60;
 buffer[503] = 8'h00;
 buffer[504] = 8'h78;
 buffer[505] = 8'hcc;
 buffer[506] = 8'h0c;
 buffer[507] = 8'h18;
 buffer[508] = 8'h30;
 buffer[509] = 8'h00;
 buffer[510] = 8'h30;
 buffer[511] = 8'h00;
 buffer[512] = 8'h7c;
 buffer[513] = 8'hc6;
 buffer[514] = 8'hde;
 buffer[515] = 8'hde;
 buffer[516] = 8'hde;
 buffer[517] = 8'hc0;
 buffer[518] = 8'h78;
 buffer[519] = 8'h00;
 buffer[520] = 8'h30;
 buffer[521] = 8'h78;
 buffer[522] = 8'hcc;
 buffer[523] = 8'hcc;
 buffer[524] = 8'hfc;
 buffer[525] = 8'hcc;
 buffer[526] = 8'hcc;
 buffer[527] = 8'h00;
 buffer[528] = 8'hfc;
 buffer[529] = 8'h66;
 buffer[530] = 8'h66;
 buffer[531] = 8'h7c;
 buffer[532] = 8'h66;
 buffer[533] = 8'h66;
 buffer[534] = 8'hfc;
 buffer[535] = 8'h00;
 buffer[536] = 8'h3c;
 buffer[537] = 8'h66;
 buffer[538] = 8'hc0;
 buffer[539] = 8'hc0;
 buffer[540] = 8'hc0;
 buffer[541] = 8'h66;
 buffer[542] = 8'h3c;
 buffer[543] = 8'h00;
 buffer[544] = 8'hf8;
 buffer[545] = 8'h6c;
 buffer[546] = 8'h66;
 buffer[547] = 8'h66;
 buffer[548] = 8'h66;
 buffer[549] = 8'h6c;
 buffer[550] = 8'hf8;
 buffer[551] = 8'h00;
 buffer[552] = 8'hfe;
 buffer[553] = 8'h62;
 buffer[554] = 8'h68;
 buffer[555] = 8'h78;
 buffer[556] = 8'h68;
 buffer[557] = 8'h62;
 buffer[558] = 8'hfe;
 buffer[559] = 8'h00;
 buffer[560] = 8'hfe;
 buffer[561] = 8'h62;
 buffer[562] = 8'h68;
 buffer[563] = 8'h78;
 buffer[564] = 8'h68;
 buffer[565] = 8'h60;
 buffer[566] = 8'hf0;
 buffer[567] = 8'h00;
 buffer[568] = 8'h3c;
 buffer[569] = 8'h66;
 buffer[570] = 8'hc0;
 buffer[571] = 8'hc0;
 buffer[572] = 8'hce;
 buffer[573] = 8'h66;
 buffer[574] = 8'h3e;
 buffer[575] = 8'h00;
 buffer[576] = 8'hcc;
 buffer[577] = 8'hcc;
 buffer[578] = 8'hcc;
 buffer[579] = 8'hfc;
 buffer[580] = 8'hcc;
 buffer[581] = 8'hcc;
 buffer[582] = 8'hcc;
 buffer[583] = 8'h00;
 buffer[584] = 8'h78;
 buffer[585] = 8'h30;
 buffer[586] = 8'h30;
 buffer[587] = 8'h30;
 buffer[588] = 8'h30;
 buffer[589] = 8'h30;
 buffer[590] = 8'h78;
 buffer[591] = 8'h00;
 buffer[592] = 8'h1e;
 buffer[593] = 8'h0c;
 buffer[594] = 8'h0c;
 buffer[595] = 8'h0c;
 buffer[596] = 8'hcc;
 buffer[597] = 8'hcc;
 buffer[598] = 8'h78;
 buffer[599] = 8'h00;
 buffer[600] = 8'he6;
 buffer[601] = 8'h66;
 buffer[602] = 8'h6c;
 buffer[603] = 8'h78;
 buffer[604] = 8'h6c;
 buffer[605] = 8'h66;
 buffer[606] = 8'he6;
 buffer[607] = 8'h00;
 buffer[608] = 8'hf0;
 buffer[609] = 8'h60;
 buffer[610] = 8'h60;
 buffer[611] = 8'h60;
 buffer[612] = 8'h62;
 buffer[613] = 8'h66;
 buffer[614] = 8'hfe;
 buffer[615] = 8'h00;
 buffer[616] = 8'hc6;
 buffer[617] = 8'hee;
 buffer[618] = 8'hfe;
 buffer[619] = 8'hfe;
 buffer[620] = 8'hd6;
 buffer[621] = 8'hc6;
 buffer[622] = 8'hc6;
 buffer[623] = 8'h00;
 buffer[624] = 8'hc6;
 buffer[625] = 8'he6;
 buffer[626] = 8'hf6;
 buffer[627] = 8'hde;
 buffer[628] = 8'hce;
 buffer[629] = 8'hc6;
 buffer[630] = 8'hc6;
 buffer[631] = 8'h00;
 buffer[632] = 8'h38;
 buffer[633] = 8'h6c;
 buffer[634] = 8'hc6;
 buffer[635] = 8'hc6;
 buffer[636] = 8'hc6;
 buffer[637] = 8'h6c;
 buffer[638] = 8'h38;
 buffer[639] = 8'h00;
 buffer[640] = 8'hfc;
 buffer[641] = 8'h66;
 buffer[642] = 8'h66;
 buffer[643] = 8'h7c;
 buffer[644] = 8'h60;
 buffer[645] = 8'h60;
 buffer[646] = 8'hf0;
 buffer[647] = 8'h00;
 buffer[648] = 8'h78;
 buffer[649] = 8'hcc;
 buffer[650] = 8'hcc;
 buffer[651] = 8'hcc;
 buffer[652] = 8'hdc;
 buffer[653] = 8'h78;
 buffer[654] = 8'h1c;
 buffer[655] = 8'h00;
 buffer[656] = 8'hfc;
 buffer[657] = 8'h66;
 buffer[658] = 8'h66;
 buffer[659] = 8'h7c;
 buffer[660] = 8'h6c;
 buffer[661] = 8'h66;
 buffer[662] = 8'he6;
 buffer[663] = 8'h00;
 buffer[664] = 8'h78;
 buffer[665] = 8'hcc;
 buffer[666] = 8'he0;
 buffer[667] = 8'h70;
 buffer[668] = 8'h1c;
 buffer[669] = 8'hcc;
 buffer[670] = 8'h78;
 buffer[671] = 8'h00;
 buffer[672] = 8'hfc;
 buffer[673] = 8'hb4;
 buffer[674] = 8'h30;
 buffer[675] = 8'h30;
 buffer[676] = 8'h30;
 buffer[677] = 8'h30;
 buffer[678] = 8'h78;
 buffer[679] = 8'h00;
 buffer[680] = 8'hcc;
 buffer[681] = 8'hcc;
 buffer[682] = 8'hcc;
 buffer[683] = 8'hcc;
 buffer[684] = 8'hcc;
 buffer[685] = 8'hcc;
 buffer[686] = 8'hfc;
 buffer[687] = 8'h00;
 buffer[688] = 8'hcc;
 buffer[689] = 8'hcc;
 buffer[690] = 8'hcc;
 buffer[691] = 8'hcc;
 buffer[692] = 8'hcc;
 buffer[693] = 8'h78;
 buffer[694] = 8'h30;
 buffer[695] = 8'h00;
 buffer[696] = 8'hc6;
 buffer[697] = 8'hc6;
 buffer[698] = 8'hc6;
 buffer[699] = 8'hd6;
 buffer[700] = 8'hfe;
 buffer[701] = 8'hee;
 buffer[702] = 8'hc6;
 buffer[703] = 8'h00;
 buffer[704] = 8'hc6;
 buffer[705] = 8'hc6;
 buffer[706] = 8'h6c;
 buffer[707] = 8'h38;
 buffer[708] = 8'h38;
 buffer[709] = 8'h6c;
 buffer[710] = 8'hc6;
 buffer[711] = 8'h00;
 buffer[712] = 8'hcc;
 buffer[713] = 8'hcc;
 buffer[714] = 8'hcc;
 buffer[715] = 8'h78;
 buffer[716] = 8'h30;
 buffer[717] = 8'h30;
 buffer[718] = 8'h78;
 buffer[719] = 8'h00;
 buffer[720] = 8'hfe;
 buffer[721] = 8'hc6;
 buffer[722] = 8'h8c;
 buffer[723] = 8'h18;
 buffer[724] = 8'h32;
 buffer[725] = 8'h66;
 buffer[726] = 8'hfe;
 buffer[727] = 8'h00;
 buffer[728] = 8'h78;
 buffer[729] = 8'h60;
 buffer[730] = 8'h60;
 buffer[731] = 8'h60;
 buffer[732] = 8'h60;
 buffer[733] = 8'h60;
 buffer[734] = 8'h78;
 buffer[735] = 8'h00;
 buffer[736] = 8'hc0;
 buffer[737] = 8'h60;
 buffer[738] = 8'h30;
 buffer[739] = 8'h18;
 buffer[740] = 8'h0c;
 buffer[741] = 8'h06;
 buffer[742] = 8'h02;
 buffer[743] = 8'h00;
 buffer[744] = 8'h78;
 buffer[745] = 8'h18;
 buffer[746] = 8'h18;
 buffer[747] = 8'h18;
 buffer[748] = 8'h18;
 buffer[749] = 8'h18;
 buffer[750] = 8'h78;
 buffer[751] = 8'h00;
 buffer[752] = 8'h10;
 buffer[753] = 8'h38;
 buffer[754] = 8'h6c;
 buffer[755] = 8'hc6;
 buffer[756] = 8'h00;
 buffer[757] = 8'h00;
 buffer[758] = 8'h00;
 buffer[759] = 8'h00;
 buffer[760] = 8'h00;
 buffer[761] = 8'h00;
 buffer[762] = 8'h00;
 buffer[763] = 8'h00;
 buffer[764] = 8'h00;
 buffer[765] = 8'h00;
 buffer[766] = 8'h00;
 buffer[767] = 8'hff;
 buffer[768] = 8'h30;
 buffer[769] = 8'h30;
 buffer[770] = 8'h18;
 buffer[771] = 8'h00;
 buffer[772] = 8'h00;
 buffer[773] = 8'h00;
 buffer[774] = 8'h00;
 buffer[775] = 8'h00;
 buffer[776] = 8'h00;
 buffer[777] = 8'h00;
 buffer[778] = 8'h78;
 buffer[779] = 8'h0c;
 buffer[780] = 8'h7c;
 buffer[781] = 8'hcc;
 buffer[782] = 8'h76;
 buffer[783] = 8'h00;
 buffer[784] = 8'he0;
 buffer[785] = 8'h60;
 buffer[786] = 8'h60;
 buffer[787] = 8'h7c;
 buffer[788] = 8'h66;
 buffer[789] = 8'h66;
 buffer[790] = 8'hdc;
 buffer[791] = 8'h00;
 buffer[792] = 8'h00;
 buffer[793] = 8'h00;
 buffer[794] = 8'h78;
 buffer[795] = 8'hcc;
 buffer[796] = 8'hc0;
 buffer[797] = 8'hcc;
 buffer[798] = 8'h78;
 buffer[799] = 8'h00;
 buffer[800] = 8'h1c;
 buffer[801] = 8'h0c;
 buffer[802] = 8'h0c;
 buffer[803] = 8'h7c;
 buffer[804] = 8'hcc;
 buffer[805] = 8'hcc;
 buffer[806] = 8'h76;
 buffer[807] = 8'h00;
 buffer[808] = 8'h00;
 buffer[809] = 8'h00;
 buffer[810] = 8'h78;
 buffer[811] = 8'hcc;
 buffer[812] = 8'hfc;
 buffer[813] = 8'hc0;
 buffer[814] = 8'h78;
 buffer[815] = 8'h00;
 buffer[816] = 8'h38;
 buffer[817] = 8'h6c;
 buffer[818] = 8'h60;
 buffer[819] = 8'hf0;
 buffer[820] = 8'h60;
 buffer[821] = 8'h60;
 buffer[822] = 8'hf0;
 buffer[823] = 8'h00;
 buffer[824] = 8'h00;
 buffer[825] = 8'h00;
 buffer[826] = 8'h76;
 buffer[827] = 8'hcc;
 buffer[828] = 8'hcc;
 buffer[829] = 8'h7c;
 buffer[830] = 8'h0c;
 buffer[831] = 8'hf8;
 buffer[832] = 8'he0;
 buffer[833] = 8'h60;
 buffer[834] = 8'h6c;
 buffer[835] = 8'h76;
 buffer[836] = 8'h66;
 buffer[837] = 8'h66;
 buffer[838] = 8'he6;
 buffer[839] = 8'h00;
 buffer[840] = 8'h30;
 buffer[841] = 8'h00;
 buffer[842] = 8'h70;
 buffer[843] = 8'h30;
 buffer[844] = 8'h30;
 buffer[845] = 8'h30;
 buffer[846] = 8'h78;
 buffer[847] = 8'h00;
 buffer[848] = 8'h0c;
 buffer[849] = 8'h00;
 buffer[850] = 8'h0c;
 buffer[851] = 8'h0c;
 buffer[852] = 8'h0c;
 buffer[853] = 8'hcc;
 buffer[854] = 8'hcc;
 buffer[855] = 8'h78;
 buffer[856] = 8'he0;
 buffer[857] = 8'h60;
 buffer[858] = 8'h66;
 buffer[859] = 8'h6c;
 buffer[860] = 8'h78;
 buffer[861] = 8'h6c;
 buffer[862] = 8'he6;
 buffer[863] = 8'h00;
 buffer[864] = 8'h70;
 buffer[865] = 8'h30;
 buffer[866] = 8'h30;
 buffer[867] = 8'h30;
 buffer[868] = 8'h30;
 buffer[869] = 8'h30;
 buffer[870] = 8'h78;
 buffer[871] = 8'h00;
 buffer[872] = 8'h00;
 buffer[873] = 8'h00;
 buffer[874] = 8'hcc;
 buffer[875] = 8'hfe;
 buffer[876] = 8'hfe;
 buffer[877] = 8'hd6;
 buffer[878] = 8'hc6;
 buffer[879] = 8'h00;
 buffer[880] = 8'h00;
 buffer[881] = 8'h00;
 buffer[882] = 8'hf8;
 buffer[883] = 8'hcc;
 buffer[884] = 8'hcc;
 buffer[885] = 8'hcc;
 buffer[886] = 8'hcc;
 buffer[887] = 8'h00;
 buffer[888] = 8'h00;
 buffer[889] = 8'h00;
 buffer[890] = 8'h78;
 buffer[891] = 8'hcc;
 buffer[892] = 8'hcc;
 buffer[893] = 8'hcc;
 buffer[894] = 8'h78;
 buffer[895] = 8'h00;
 buffer[896] = 8'h00;
 buffer[897] = 8'h00;
 buffer[898] = 8'hdc;
 buffer[899] = 8'h66;
 buffer[900] = 8'h66;
 buffer[901] = 8'h7c;
 buffer[902] = 8'h60;
 buffer[903] = 8'hf0;
 buffer[904] = 8'h00;
 buffer[905] = 8'h00;
 buffer[906] = 8'h76;
 buffer[907] = 8'hcc;
 buffer[908] = 8'hcc;
 buffer[909] = 8'h7c;
 buffer[910] = 8'h0c;
 buffer[911] = 8'h1e;
 buffer[912] = 8'h00;
 buffer[913] = 8'h00;
 buffer[914] = 8'hdc;
 buffer[915] = 8'h76;
 buffer[916] = 8'h66;
 buffer[917] = 8'h60;
 buffer[918] = 8'hf0;
 buffer[919] = 8'h00;
 buffer[920] = 8'h00;
 buffer[921] = 8'h00;
 buffer[922] = 8'h7c;
 buffer[923] = 8'hc0;
 buffer[924] = 8'h78;
 buffer[925] = 8'h0c;
 buffer[926] = 8'hf8;
 buffer[927] = 8'h00;
 buffer[928] = 8'h10;
 buffer[929] = 8'h30;
 buffer[930] = 8'h7c;
 buffer[931] = 8'h30;
 buffer[932] = 8'h30;
 buffer[933] = 8'h34;
 buffer[934] = 8'h18;
 buffer[935] = 8'h00;
 buffer[936] = 8'h00;
 buffer[937] = 8'h00;
 buffer[938] = 8'hcc;
 buffer[939] = 8'hcc;
 buffer[940] = 8'hcc;
 buffer[941] = 8'hcc;
 buffer[942] = 8'h76;
 buffer[943] = 8'h00;
 buffer[944] = 8'h00;
 buffer[945] = 8'h00;
 buffer[946] = 8'hcc;
 buffer[947] = 8'hcc;
 buffer[948] = 8'hcc;
 buffer[949] = 8'h78;
 buffer[950] = 8'h30;
 buffer[951] = 8'h00;
 buffer[952] = 8'h00;
 buffer[953] = 8'h00;
 buffer[954] = 8'hc6;
 buffer[955] = 8'hd6;
 buffer[956] = 8'hfe;
 buffer[957] = 8'hfe;
 buffer[958] = 8'h6c;
 buffer[959] = 8'h00;
 buffer[960] = 8'h00;
 buffer[961] = 8'h00;
 buffer[962] = 8'hc6;
 buffer[963] = 8'h6c;
 buffer[964] = 8'h38;
 buffer[965] = 8'h6c;
 buffer[966] = 8'hc6;
 buffer[967] = 8'h00;
 buffer[968] = 8'h00;
 buffer[969] = 8'h00;
 buffer[970] = 8'hcc;
 buffer[971] = 8'hcc;
 buffer[972] = 8'hcc;
 buffer[973] = 8'h7c;
 buffer[974] = 8'h0c;
 buffer[975] = 8'hf8;
 buffer[976] = 8'h00;
 buffer[977] = 8'h00;
 buffer[978] = 8'hfc;
 buffer[979] = 8'h98;
 buffer[980] = 8'h30;
 buffer[981] = 8'h64;
 buffer[982] = 8'hfc;
 buffer[983] = 8'h00;
 buffer[984] = 8'h1c;
 buffer[985] = 8'h30;
 buffer[986] = 8'h30;
 buffer[987] = 8'he0;
 buffer[988] = 8'h30;
 buffer[989] = 8'h30;
 buffer[990] = 8'h1c;
 buffer[991] = 8'h00;
 buffer[992] = 8'h18;
 buffer[993] = 8'h18;
 buffer[994] = 8'h18;
 buffer[995] = 8'h00;
 buffer[996] = 8'h18;
 buffer[997] = 8'h18;
 buffer[998] = 8'h18;
 buffer[999] = 8'h00;
 buffer[1000] = 8'he0;
 buffer[1001] = 8'h30;
 buffer[1002] = 8'h30;
 buffer[1003] = 8'h1c;
 buffer[1004] = 8'h30;
 buffer[1005] = 8'h30;
 buffer[1006] = 8'he0;
 buffer[1007] = 8'h00;
 buffer[1008] = 8'h76;
 buffer[1009] = 8'hdc;
 buffer[1010] = 8'h00;
 buffer[1011] = 8'h00;
 buffer[1012] = 8'h00;
 buffer[1013] = 8'h00;
 buffer[1014] = 8'h00;
 buffer[1015] = 8'h00;
 buffer[1016] = 8'h00;
 buffer[1017] = 8'h10;
 buffer[1018] = 8'h38;
 buffer[1019] = 8'h6c;
 buffer[1020] = 8'hc6;
 buffer[1021] = 8'hc6;
 buffer[1022] = 8'hfe;
 buffer[1023] = 8'h00;
 buffer[1024] = 8'h78;
 buffer[1025] = 8'hcc;
 buffer[1026] = 8'hc0;
 buffer[1027] = 8'hcc;
 buffer[1028] = 8'h78;
 buffer[1029] = 8'h18;
 buffer[1030] = 8'h0c;
 buffer[1031] = 8'h78;
 buffer[1032] = 8'h00;
 buffer[1033] = 8'hcc;
 buffer[1034] = 8'h00;
 buffer[1035] = 8'hcc;
 buffer[1036] = 8'hcc;
 buffer[1037] = 8'hcc;
 buffer[1038] = 8'h7e;
 buffer[1039] = 8'h00;
 buffer[1040] = 8'h1c;
 buffer[1041] = 8'h00;
 buffer[1042] = 8'h78;
 buffer[1043] = 8'hcc;
 buffer[1044] = 8'hfc;
 buffer[1045] = 8'hc0;
 buffer[1046] = 8'h78;
 buffer[1047] = 8'h00;
 buffer[1048] = 8'h7e;
 buffer[1049] = 8'hc3;
 buffer[1050] = 8'h3c;
 buffer[1051] = 8'h06;
 buffer[1052] = 8'h3e;
 buffer[1053] = 8'h66;
 buffer[1054] = 8'h3f;
 buffer[1055] = 8'h00;
 buffer[1056] = 8'hcc;
 buffer[1057] = 8'h00;
 buffer[1058] = 8'h78;
 buffer[1059] = 8'h0c;
 buffer[1060] = 8'h7c;
 buffer[1061] = 8'hcc;
 buffer[1062] = 8'h7e;
 buffer[1063] = 8'h00;
 buffer[1064] = 8'he0;
 buffer[1065] = 8'h00;
 buffer[1066] = 8'h78;
 buffer[1067] = 8'h0c;
 buffer[1068] = 8'h7c;
 buffer[1069] = 8'hcc;
 buffer[1070] = 8'h7e;
 buffer[1071] = 8'h00;
 buffer[1072] = 8'h30;
 buffer[1073] = 8'h30;
 buffer[1074] = 8'h78;
 buffer[1075] = 8'h0c;
 buffer[1076] = 8'h7c;
 buffer[1077] = 8'hcc;
 buffer[1078] = 8'h7e;
 buffer[1079] = 8'h00;
 buffer[1080] = 8'h00;
 buffer[1081] = 8'h00;
 buffer[1082] = 8'h78;
 buffer[1083] = 8'hc0;
 buffer[1084] = 8'hc0;
 buffer[1085] = 8'h78;
 buffer[1086] = 8'h0c;
 buffer[1087] = 8'h38;
 buffer[1088] = 8'h7e;
 buffer[1089] = 8'hc3;
 buffer[1090] = 8'h3c;
 buffer[1091] = 8'h66;
 buffer[1092] = 8'h7e;
 buffer[1093] = 8'h60;
 buffer[1094] = 8'h3c;
 buffer[1095] = 8'h00;
 buffer[1096] = 8'hcc;
 buffer[1097] = 8'h00;
 buffer[1098] = 8'h78;
 buffer[1099] = 8'hcc;
 buffer[1100] = 8'hfc;
 buffer[1101] = 8'hc0;
 buffer[1102] = 8'h78;
 buffer[1103] = 8'h00;
 buffer[1104] = 8'he0;
 buffer[1105] = 8'h00;
 buffer[1106] = 8'h78;
 buffer[1107] = 8'hcc;
 buffer[1108] = 8'hfc;
 buffer[1109] = 8'hc0;
 buffer[1110] = 8'h78;
 buffer[1111] = 8'h00;
 buffer[1112] = 8'hcc;
 buffer[1113] = 8'h00;
 buffer[1114] = 8'h70;
 buffer[1115] = 8'h30;
 buffer[1116] = 8'h30;
 buffer[1117] = 8'h30;
 buffer[1118] = 8'h78;
 buffer[1119] = 8'h00;
 buffer[1120] = 8'h7c;
 buffer[1121] = 8'hc6;
 buffer[1122] = 8'h38;
 buffer[1123] = 8'h18;
 buffer[1124] = 8'h18;
 buffer[1125] = 8'h18;
 buffer[1126] = 8'h3c;
 buffer[1127] = 8'h00;
 buffer[1128] = 8'he0;
 buffer[1129] = 8'h00;
 buffer[1130] = 8'h70;
 buffer[1131] = 8'h30;
 buffer[1132] = 8'h30;
 buffer[1133] = 8'h30;
 buffer[1134] = 8'h78;
 buffer[1135] = 8'h00;
 buffer[1136] = 8'hc6;
 buffer[1137] = 8'h38;
 buffer[1138] = 8'h6c;
 buffer[1139] = 8'hc6;
 buffer[1140] = 8'hfe;
 buffer[1141] = 8'hc6;
 buffer[1142] = 8'hc6;
 buffer[1143] = 8'h00;
 buffer[1144] = 8'h30;
 buffer[1145] = 8'h30;
 buffer[1146] = 8'h00;
 buffer[1147] = 8'h78;
 buffer[1148] = 8'hcc;
 buffer[1149] = 8'hfc;
 buffer[1150] = 8'hcc;
 buffer[1151] = 8'h00;
 buffer[1152] = 8'h1c;
 buffer[1153] = 8'h00;
 buffer[1154] = 8'hfc;
 buffer[1155] = 8'h60;
 buffer[1156] = 8'h78;
 buffer[1157] = 8'h60;
 buffer[1158] = 8'hfc;
 buffer[1159] = 8'h00;
 buffer[1160] = 8'h00;
 buffer[1161] = 8'h00;
 buffer[1162] = 8'h7f;
 buffer[1163] = 8'h0c;
 buffer[1164] = 8'h7f;
 buffer[1165] = 8'hcc;
 buffer[1166] = 8'h7f;
 buffer[1167] = 8'h00;
 buffer[1168] = 8'h3e;
 buffer[1169] = 8'h6c;
 buffer[1170] = 8'hcc;
 buffer[1171] = 8'hfe;
 buffer[1172] = 8'hcc;
 buffer[1173] = 8'hcc;
 buffer[1174] = 8'hce;
 buffer[1175] = 8'h00;
 buffer[1176] = 8'h78;
 buffer[1177] = 8'hcc;
 buffer[1178] = 8'h00;
 buffer[1179] = 8'h78;
 buffer[1180] = 8'hcc;
 buffer[1181] = 8'hcc;
 buffer[1182] = 8'h78;
 buffer[1183] = 8'h00;
 buffer[1184] = 8'h00;
 buffer[1185] = 8'hcc;
 buffer[1186] = 8'h00;
 buffer[1187] = 8'h78;
 buffer[1188] = 8'hcc;
 buffer[1189] = 8'hcc;
 buffer[1190] = 8'h78;
 buffer[1191] = 8'h00;
 buffer[1192] = 8'h00;
 buffer[1193] = 8'he0;
 buffer[1194] = 8'h00;
 buffer[1195] = 8'h78;
 buffer[1196] = 8'hcc;
 buffer[1197] = 8'hcc;
 buffer[1198] = 8'h78;
 buffer[1199] = 8'h00;
 buffer[1200] = 8'h78;
 buffer[1201] = 8'hcc;
 buffer[1202] = 8'h00;
 buffer[1203] = 8'hcc;
 buffer[1204] = 8'hcc;
 buffer[1205] = 8'hcc;
 buffer[1206] = 8'h7e;
 buffer[1207] = 8'h00;
 buffer[1208] = 8'h00;
 buffer[1209] = 8'he0;
 buffer[1210] = 8'h00;
 buffer[1211] = 8'hcc;
 buffer[1212] = 8'hcc;
 buffer[1213] = 8'hcc;
 buffer[1214] = 8'h7e;
 buffer[1215] = 8'h00;
 buffer[1216] = 8'h00;
 buffer[1217] = 8'hcc;
 buffer[1218] = 8'h00;
 buffer[1219] = 8'hcc;
 buffer[1220] = 8'hcc;
 buffer[1221] = 8'h7c;
 buffer[1222] = 8'h0c;
 buffer[1223] = 8'hf8;
 buffer[1224] = 8'hc3;
 buffer[1225] = 8'h18;
 buffer[1226] = 8'h3c;
 buffer[1227] = 8'h66;
 buffer[1228] = 8'h66;
 buffer[1229] = 8'h3c;
 buffer[1230] = 8'h18;
 buffer[1231] = 8'h00;
 buffer[1232] = 8'hcc;
 buffer[1233] = 8'h00;
 buffer[1234] = 8'hcc;
 buffer[1235] = 8'hcc;
 buffer[1236] = 8'hcc;
 buffer[1237] = 8'hcc;
 buffer[1238] = 8'h78;
 buffer[1239] = 8'h00;
 buffer[1240] = 8'h18;
 buffer[1241] = 8'h18;
 buffer[1242] = 8'h7e;
 buffer[1243] = 8'hc0;
 buffer[1244] = 8'hc0;
 buffer[1245] = 8'h7e;
 buffer[1246] = 8'h18;
 buffer[1247] = 8'h18;
 buffer[1248] = 8'h38;
 buffer[1249] = 8'h6c;
 buffer[1250] = 8'h64;
 buffer[1251] = 8'hf0;
 buffer[1252] = 8'h60;
 buffer[1253] = 8'he6;
 buffer[1254] = 8'hfc;
 buffer[1255] = 8'h00;
 buffer[1256] = 8'hcc;
 buffer[1257] = 8'hcc;
 buffer[1258] = 8'h78;
 buffer[1259] = 8'hfc;
 buffer[1260] = 8'h30;
 buffer[1261] = 8'hfc;
 buffer[1262] = 8'h30;
 buffer[1263] = 8'h30;
 buffer[1264] = 8'hf8;
 buffer[1265] = 8'hcc;
 buffer[1266] = 8'hcc;
 buffer[1267] = 8'hfa;
 buffer[1268] = 8'hc6;
 buffer[1269] = 8'hcf;
 buffer[1270] = 8'hc6;
 buffer[1271] = 8'hc7;
 buffer[1272] = 8'h0e;
 buffer[1273] = 8'h1b;
 buffer[1274] = 8'h18;
 buffer[1275] = 8'h3c;
 buffer[1276] = 8'h18;
 buffer[1277] = 8'h18;
 buffer[1278] = 8'hd8;
 buffer[1279] = 8'h70;
 buffer[1280] = 8'h1c;
 buffer[1281] = 8'h00;
 buffer[1282] = 8'h78;
 buffer[1283] = 8'h0c;
 buffer[1284] = 8'h7c;
 buffer[1285] = 8'hcc;
 buffer[1286] = 8'h7e;
 buffer[1287] = 8'h00;
 buffer[1288] = 8'h38;
 buffer[1289] = 8'h00;
 buffer[1290] = 8'h70;
 buffer[1291] = 8'h30;
 buffer[1292] = 8'h30;
 buffer[1293] = 8'h30;
 buffer[1294] = 8'h78;
 buffer[1295] = 8'h00;
 buffer[1296] = 8'h00;
 buffer[1297] = 8'h1c;
 buffer[1298] = 8'h00;
 buffer[1299] = 8'h78;
 buffer[1300] = 8'hcc;
 buffer[1301] = 8'hcc;
 buffer[1302] = 8'h78;
 buffer[1303] = 8'h00;
 buffer[1304] = 8'h00;
 buffer[1305] = 8'h1c;
 buffer[1306] = 8'h00;
 buffer[1307] = 8'hcc;
 buffer[1308] = 8'hcc;
 buffer[1309] = 8'hcc;
 buffer[1310] = 8'h7e;
 buffer[1311] = 8'h00;
 buffer[1312] = 8'h00;
 buffer[1313] = 8'hf8;
 buffer[1314] = 8'h00;
 buffer[1315] = 8'hf8;
 buffer[1316] = 8'hcc;
 buffer[1317] = 8'hcc;
 buffer[1318] = 8'hcc;
 buffer[1319] = 8'h00;
 buffer[1320] = 8'hfc;
 buffer[1321] = 8'h00;
 buffer[1322] = 8'hcc;
 buffer[1323] = 8'hec;
 buffer[1324] = 8'hfc;
 buffer[1325] = 8'hdc;
 buffer[1326] = 8'hcc;
 buffer[1327] = 8'h00;
 buffer[1328] = 8'h3c;
 buffer[1329] = 8'h6c;
 buffer[1330] = 8'h6c;
 buffer[1331] = 8'h3e;
 buffer[1332] = 8'h00;
 buffer[1333] = 8'h7e;
 buffer[1334] = 8'h00;
 buffer[1335] = 8'h00;
 buffer[1336] = 8'h38;
 buffer[1337] = 8'h6c;
 buffer[1338] = 8'h6c;
 buffer[1339] = 8'h38;
 buffer[1340] = 8'h00;
 buffer[1341] = 8'h7c;
 buffer[1342] = 8'h00;
 buffer[1343] = 8'h00;
 buffer[1344] = 8'h30;
 buffer[1345] = 8'h00;
 buffer[1346] = 8'h30;
 buffer[1347] = 8'h60;
 buffer[1348] = 8'hc0;
 buffer[1349] = 8'hcc;
 buffer[1350] = 8'h78;
 buffer[1351] = 8'h00;
 buffer[1352] = 8'h00;
 buffer[1353] = 8'h00;
 buffer[1354] = 8'h00;
 buffer[1355] = 8'hfc;
 buffer[1356] = 8'hc0;
 buffer[1357] = 8'hc0;
 buffer[1358] = 8'h00;
 buffer[1359] = 8'h00;
 buffer[1360] = 8'h00;
 buffer[1361] = 8'h00;
 buffer[1362] = 8'h00;
 buffer[1363] = 8'hfc;
 buffer[1364] = 8'h0c;
 buffer[1365] = 8'h0c;
 buffer[1366] = 8'h00;
 buffer[1367] = 8'h00;
 buffer[1368] = 8'hc3;
 buffer[1369] = 8'hc6;
 buffer[1370] = 8'hcc;
 buffer[1371] = 8'hde;
 buffer[1372] = 8'h33;
 buffer[1373] = 8'h66;
 buffer[1374] = 8'hcc;
 buffer[1375] = 8'h0f;
 buffer[1376] = 8'hc3;
 buffer[1377] = 8'hc6;
 buffer[1378] = 8'hcc;
 buffer[1379] = 8'hdb;
 buffer[1380] = 8'h37;
 buffer[1381] = 8'h6f;
 buffer[1382] = 8'hcf;
 buffer[1383] = 8'h03;
 buffer[1384] = 8'h18;
 buffer[1385] = 8'h18;
 buffer[1386] = 8'h00;
 buffer[1387] = 8'h18;
 buffer[1388] = 8'h18;
 buffer[1389] = 8'h18;
 buffer[1390] = 8'h18;
 buffer[1391] = 8'h00;
 buffer[1392] = 8'h00;
 buffer[1393] = 8'h33;
 buffer[1394] = 8'h66;
 buffer[1395] = 8'hcc;
 buffer[1396] = 8'h66;
 buffer[1397] = 8'h33;
 buffer[1398] = 8'h00;
 buffer[1399] = 8'h00;
 buffer[1400] = 8'h00;
 buffer[1401] = 8'hcc;
 buffer[1402] = 8'h66;
 buffer[1403] = 8'h33;
 buffer[1404] = 8'h66;
 buffer[1405] = 8'hcc;
 buffer[1406] = 8'h00;
 buffer[1407] = 8'h00;
 buffer[1408] = 8'h22;
 buffer[1409] = 8'h88;
 buffer[1410] = 8'h22;
 buffer[1411] = 8'h88;
 buffer[1412] = 8'h22;
 buffer[1413] = 8'h88;
 buffer[1414] = 8'h22;
 buffer[1415] = 8'h88;
 buffer[1416] = 8'h55;
 buffer[1417] = 8'haa;
 buffer[1418] = 8'h55;
 buffer[1419] = 8'haa;
 buffer[1420] = 8'h55;
 buffer[1421] = 8'haa;
 buffer[1422] = 8'h55;
 buffer[1423] = 8'haa;
 buffer[1424] = 8'hdb;
 buffer[1425] = 8'h77;
 buffer[1426] = 8'hdb;
 buffer[1427] = 8'hee;
 buffer[1428] = 8'hdb;
 buffer[1429] = 8'h77;
 buffer[1430] = 8'hdb;
 buffer[1431] = 8'hee;
 buffer[1432] = 8'h18;
 buffer[1433] = 8'h18;
 buffer[1434] = 8'h18;
 buffer[1435] = 8'h18;
 buffer[1436] = 8'h18;
 buffer[1437] = 8'h18;
 buffer[1438] = 8'h18;
 buffer[1439] = 8'h18;
 buffer[1440] = 8'h18;
 buffer[1441] = 8'h18;
 buffer[1442] = 8'h18;
 buffer[1443] = 8'h18;
 buffer[1444] = 8'hf8;
 buffer[1445] = 8'h18;
 buffer[1446] = 8'h18;
 buffer[1447] = 8'h18;
 buffer[1448] = 8'h18;
 buffer[1449] = 8'h18;
 buffer[1450] = 8'hf8;
 buffer[1451] = 8'h18;
 buffer[1452] = 8'hf8;
 buffer[1453] = 8'h18;
 buffer[1454] = 8'h18;
 buffer[1455] = 8'h18;
 buffer[1456] = 8'h36;
 buffer[1457] = 8'h36;
 buffer[1458] = 8'h36;
 buffer[1459] = 8'h36;
 buffer[1460] = 8'hf6;
 buffer[1461] = 8'h36;
 buffer[1462] = 8'h36;
 buffer[1463] = 8'h36;
 buffer[1464] = 8'h00;
 buffer[1465] = 8'h00;
 buffer[1466] = 8'h00;
 buffer[1467] = 8'h00;
 buffer[1468] = 8'hfe;
 buffer[1469] = 8'h36;
 buffer[1470] = 8'h36;
 buffer[1471] = 8'h36;
 buffer[1472] = 8'h00;
 buffer[1473] = 8'h00;
 buffer[1474] = 8'hf8;
 buffer[1475] = 8'h18;
 buffer[1476] = 8'hf8;
 buffer[1477] = 8'h18;
 buffer[1478] = 8'h18;
 buffer[1479] = 8'h18;
 buffer[1480] = 8'h36;
 buffer[1481] = 8'h36;
 buffer[1482] = 8'hf6;
 buffer[1483] = 8'h06;
 buffer[1484] = 8'hf6;
 buffer[1485] = 8'h36;
 buffer[1486] = 8'h36;
 buffer[1487] = 8'h36;
 buffer[1488] = 8'h36;
 buffer[1489] = 8'h36;
 buffer[1490] = 8'h36;
 buffer[1491] = 8'h36;
 buffer[1492] = 8'h36;
 buffer[1493] = 8'h36;
 buffer[1494] = 8'h36;
 buffer[1495] = 8'h36;
 buffer[1496] = 8'h00;
 buffer[1497] = 8'h00;
 buffer[1498] = 8'hfe;
 buffer[1499] = 8'h06;
 buffer[1500] = 8'hf6;
 buffer[1501] = 8'h36;
 buffer[1502] = 8'h36;
 buffer[1503] = 8'h36;
 buffer[1504] = 8'h36;
 buffer[1505] = 8'h36;
 buffer[1506] = 8'hf6;
 buffer[1507] = 8'h06;
 buffer[1508] = 8'hfe;
 buffer[1509] = 8'h00;
 buffer[1510] = 8'h00;
 buffer[1511] = 8'h00;
 buffer[1512] = 8'h36;
 buffer[1513] = 8'h36;
 buffer[1514] = 8'h36;
 buffer[1515] = 8'h36;
 buffer[1516] = 8'hfe;
 buffer[1517] = 8'h00;
 buffer[1518] = 8'h00;
 buffer[1519] = 8'h00;
 buffer[1520] = 8'h18;
 buffer[1521] = 8'h18;
 buffer[1522] = 8'hf8;
 buffer[1523] = 8'h18;
 buffer[1524] = 8'hf8;
 buffer[1525] = 8'h00;
 buffer[1526] = 8'h00;
 buffer[1527] = 8'h00;
 buffer[1528] = 8'h00;
 buffer[1529] = 8'h00;
 buffer[1530] = 8'h00;
 buffer[1531] = 8'h00;
 buffer[1532] = 8'hf8;
 buffer[1533] = 8'h18;
 buffer[1534] = 8'h18;
 buffer[1535] = 8'h18;
 buffer[1536] = 8'h18;
 buffer[1537] = 8'h18;
 buffer[1538] = 8'h18;
 buffer[1539] = 8'h18;
 buffer[1540] = 8'h1f;
 buffer[1541] = 8'h00;
 buffer[1542] = 8'h00;
 buffer[1543] = 8'h00;
 buffer[1544] = 8'h18;
 buffer[1545] = 8'h18;
 buffer[1546] = 8'h18;
 buffer[1547] = 8'h18;
 buffer[1548] = 8'hff;
 buffer[1549] = 8'h00;
 buffer[1550] = 8'h00;
 buffer[1551] = 8'h00;
 buffer[1552] = 8'h00;
 buffer[1553] = 8'h00;
 buffer[1554] = 8'h00;
 buffer[1555] = 8'h00;
 buffer[1556] = 8'hff;
 buffer[1557] = 8'h18;
 buffer[1558] = 8'h18;
 buffer[1559] = 8'h18;
 buffer[1560] = 8'h18;
 buffer[1561] = 8'h18;
 buffer[1562] = 8'h18;
 buffer[1563] = 8'h18;
 buffer[1564] = 8'h1f;
 buffer[1565] = 8'h18;
 buffer[1566] = 8'h18;
 buffer[1567] = 8'h18;
 buffer[1568] = 8'h00;
 buffer[1569] = 8'h00;
 buffer[1570] = 8'h00;
 buffer[1571] = 8'h00;
 buffer[1572] = 8'hff;
 buffer[1573] = 8'h00;
 buffer[1574] = 8'h00;
 buffer[1575] = 8'h00;
 buffer[1576] = 8'h18;
 buffer[1577] = 8'h18;
 buffer[1578] = 8'h18;
 buffer[1579] = 8'h18;
 buffer[1580] = 8'hff;
 buffer[1581] = 8'h18;
 buffer[1582] = 8'h18;
 buffer[1583] = 8'h18;
 buffer[1584] = 8'h18;
 buffer[1585] = 8'h18;
 buffer[1586] = 8'h1f;
 buffer[1587] = 8'h18;
 buffer[1588] = 8'h1f;
 buffer[1589] = 8'h18;
 buffer[1590] = 8'h18;
 buffer[1591] = 8'h18;
 buffer[1592] = 8'h36;
 buffer[1593] = 8'h36;
 buffer[1594] = 8'h36;
 buffer[1595] = 8'h36;
 buffer[1596] = 8'h37;
 buffer[1597] = 8'h36;
 buffer[1598] = 8'h36;
 buffer[1599] = 8'h36;
 buffer[1600] = 8'h36;
 buffer[1601] = 8'h36;
 buffer[1602] = 8'h37;
 buffer[1603] = 8'h30;
 buffer[1604] = 8'h3f;
 buffer[1605] = 8'h00;
 buffer[1606] = 8'h00;
 buffer[1607] = 8'h00;
 buffer[1608] = 8'h00;
 buffer[1609] = 8'h00;
 buffer[1610] = 8'h3f;
 buffer[1611] = 8'h30;
 buffer[1612] = 8'h37;
 buffer[1613] = 8'h36;
 buffer[1614] = 8'h36;
 buffer[1615] = 8'h36;
 buffer[1616] = 8'h36;
 buffer[1617] = 8'h36;
 buffer[1618] = 8'hf7;
 buffer[1619] = 8'h00;
 buffer[1620] = 8'hff;
 buffer[1621] = 8'h00;
 buffer[1622] = 8'h00;
 buffer[1623] = 8'h00;
 buffer[1624] = 8'h00;
 buffer[1625] = 8'h00;
 buffer[1626] = 8'hff;
 buffer[1627] = 8'h00;
 buffer[1628] = 8'hf7;
 buffer[1629] = 8'h36;
 buffer[1630] = 8'h36;
 buffer[1631] = 8'h36;
 buffer[1632] = 8'h36;
 buffer[1633] = 8'h36;
 buffer[1634] = 8'h37;
 buffer[1635] = 8'h30;
 buffer[1636] = 8'h37;
 buffer[1637] = 8'h36;
 buffer[1638] = 8'h36;
 buffer[1639] = 8'h36;
 buffer[1640] = 8'h00;
 buffer[1641] = 8'h00;
 buffer[1642] = 8'hff;
 buffer[1643] = 8'h00;
 buffer[1644] = 8'hff;
 buffer[1645] = 8'h00;
 buffer[1646] = 8'h00;
 buffer[1647] = 8'h00;
 buffer[1648] = 8'h36;
 buffer[1649] = 8'h36;
 buffer[1650] = 8'hf7;
 buffer[1651] = 8'h00;
 buffer[1652] = 8'hf7;
 buffer[1653] = 8'h36;
 buffer[1654] = 8'h36;
 buffer[1655] = 8'h36;
 buffer[1656] = 8'h18;
 buffer[1657] = 8'h18;
 buffer[1658] = 8'hff;
 buffer[1659] = 8'h00;
 buffer[1660] = 8'hff;
 buffer[1661] = 8'h00;
 buffer[1662] = 8'h00;
 buffer[1663] = 8'h00;
 buffer[1664] = 8'h36;
 buffer[1665] = 8'h36;
 buffer[1666] = 8'h36;
 buffer[1667] = 8'h36;
 buffer[1668] = 8'hff;
 buffer[1669] = 8'h00;
 buffer[1670] = 8'h00;
 buffer[1671] = 8'h00;
 buffer[1672] = 8'h00;
 buffer[1673] = 8'h00;
 buffer[1674] = 8'hff;
 buffer[1675] = 8'h00;
 buffer[1676] = 8'hff;
 buffer[1677] = 8'h18;
 buffer[1678] = 8'h18;
 buffer[1679] = 8'h18;
 buffer[1680] = 8'h00;
 buffer[1681] = 8'h00;
 buffer[1682] = 8'h00;
 buffer[1683] = 8'h00;
 buffer[1684] = 8'hff;
 buffer[1685] = 8'h36;
 buffer[1686] = 8'h36;
 buffer[1687] = 8'h36;
 buffer[1688] = 8'h36;
 buffer[1689] = 8'h36;
 buffer[1690] = 8'h36;
 buffer[1691] = 8'h36;
 buffer[1692] = 8'h3f;
 buffer[1693] = 8'h00;
 buffer[1694] = 8'h00;
 buffer[1695] = 8'h00;
 buffer[1696] = 8'h18;
 buffer[1697] = 8'h18;
 buffer[1698] = 8'h1f;
 buffer[1699] = 8'h18;
 buffer[1700] = 8'h1f;
 buffer[1701] = 8'h00;
 buffer[1702] = 8'h00;
 buffer[1703] = 8'h00;
 buffer[1704] = 8'h00;
 buffer[1705] = 8'h00;
 buffer[1706] = 8'h1f;
 buffer[1707] = 8'h18;
 buffer[1708] = 8'h1f;
 buffer[1709] = 8'h18;
 buffer[1710] = 8'h18;
 buffer[1711] = 8'h18;
 buffer[1712] = 8'h00;
 buffer[1713] = 8'h00;
 buffer[1714] = 8'h00;
 buffer[1715] = 8'h00;
 buffer[1716] = 8'h3f;
 buffer[1717] = 8'h36;
 buffer[1718] = 8'h36;
 buffer[1719] = 8'h36;
 buffer[1720] = 8'h36;
 buffer[1721] = 8'h36;
 buffer[1722] = 8'h36;
 buffer[1723] = 8'h36;
 buffer[1724] = 8'hff;
 buffer[1725] = 8'h36;
 buffer[1726] = 8'h36;
 buffer[1727] = 8'h36;
 buffer[1728] = 8'h18;
 buffer[1729] = 8'h18;
 buffer[1730] = 8'hff;
 buffer[1731] = 8'h18;
 buffer[1732] = 8'hff;
 buffer[1733] = 8'h18;
 buffer[1734] = 8'h18;
 buffer[1735] = 8'h18;
 buffer[1736] = 8'h18;
 buffer[1737] = 8'h18;
 buffer[1738] = 8'h18;
 buffer[1739] = 8'h18;
 buffer[1740] = 8'hf8;
 buffer[1741] = 8'h00;
 buffer[1742] = 8'h00;
 buffer[1743] = 8'h00;
 buffer[1744] = 8'h00;
 buffer[1745] = 8'h00;
 buffer[1746] = 8'h00;
 buffer[1747] = 8'h00;
 buffer[1748] = 8'h1f;
 buffer[1749] = 8'h18;
 buffer[1750] = 8'h18;
 buffer[1751] = 8'h18;
 buffer[1752] = 8'hff;
 buffer[1753] = 8'hff;
 buffer[1754] = 8'hff;
 buffer[1755] = 8'hff;
 buffer[1756] = 8'hff;
 buffer[1757] = 8'hff;
 buffer[1758] = 8'hff;
 buffer[1759] = 8'hff;
 buffer[1760] = 8'h00;
 buffer[1761] = 8'h00;
 buffer[1762] = 8'h00;
 buffer[1763] = 8'h00;
 buffer[1764] = 8'hff;
 buffer[1765] = 8'hff;
 buffer[1766] = 8'hff;
 buffer[1767] = 8'hff;
 buffer[1768] = 8'hf0;
 buffer[1769] = 8'hf0;
 buffer[1770] = 8'hf0;
 buffer[1771] = 8'hf0;
 buffer[1772] = 8'hf0;
 buffer[1773] = 8'hf0;
 buffer[1774] = 8'hf0;
 buffer[1775] = 8'hf0;
 buffer[1776] = 8'h0f;
 buffer[1777] = 8'h0f;
 buffer[1778] = 8'h0f;
 buffer[1779] = 8'h0f;
 buffer[1780] = 8'h0f;
 buffer[1781] = 8'h0f;
 buffer[1782] = 8'h0f;
 buffer[1783] = 8'h0f;
 buffer[1784] = 8'hff;
 buffer[1785] = 8'hff;
 buffer[1786] = 8'hff;
 buffer[1787] = 8'hff;
 buffer[1788] = 8'h00;
 buffer[1789] = 8'h00;
 buffer[1790] = 8'h00;
 buffer[1791] = 8'h00;
 buffer[1792] = 8'h00;
 buffer[1793] = 8'h00;
 buffer[1794] = 8'h76;
 buffer[1795] = 8'hdc;
 buffer[1796] = 8'hc8;
 buffer[1797] = 8'hdc;
 buffer[1798] = 8'h76;
 buffer[1799] = 8'h00;
 buffer[1800] = 8'h00;
 buffer[1801] = 8'h78;
 buffer[1802] = 8'hcc;
 buffer[1803] = 8'hf8;
 buffer[1804] = 8'hcc;
 buffer[1805] = 8'hf8;
 buffer[1806] = 8'hc0;
 buffer[1807] = 8'hc0;
 buffer[1808] = 8'h00;
 buffer[1809] = 8'hfc;
 buffer[1810] = 8'hcc;
 buffer[1811] = 8'hc0;
 buffer[1812] = 8'hc0;
 buffer[1813] = 8'hc0;
 buffer[1814] = 8'hc0;
 buffer[1815] = 8'h00;
 buffer[1816] = 8'h00;
 buffer[1817] = 8'hfe;
 buffer[1818] = 8'h6c;
 buffer[1819] = 8'h6c;
 buffer[1820] = 8'h6c;
 buffer[1821] = 8'h6c;
 buffer[1822] = 8'h6c;
 buffer[1823] = 8'h00;
 buffer[1824] = 8'hfc;
 buffer[1825] = 8'hcc;
 buffer[1826] = 8'h60;
 buffer[1827] = 8'h30;
 buffer[1828] = 8'h60;
 buffer[1829] = 8'hcc;
 buffer[1830] = 8'hfc;
 buffer[1831] = 8'h00;
 buffer[1832] = 8'h00;
 buffer[1833] = 8'h00;
 buffer[1834] = 8'h7e;
 buffer[1835] = 8'hd8;
 buffer[1836] = 8'hd8;
 buffer[1837] = 8'hd8;
 buffer[1838] = 8'h70;
 buffer[1839] = 8'h00;
 buffer[1840] = 8'h00;
 buffer[1841] = 8'h66;
 buffer[1842] = 8'h66;
 buffer[1843] = 8'h66;
 buffer[1844] = 8'h66;
 buffer[1845] = 8'h7c;
 buffer[1846] = 8'h60;
 buffer[1847] = 8'hc0;
 buffer[1848] = 8'h00;
 buffer[1849] = 8'h76;
 buffer[1850] = 8'hdc;
 buffer[1851] = 8'h18;
 buffer[1852] = 8'h18;
 buffer[1853] = 8'h18;
 buffer[1854] = 8'h18;
 buffer[1855] = 8'h00;
 buffer[1856] = 8'hfc;
 buffer[1857] = 8'h30;
 buffer[1858] = 8'h78;
 buffer[1859] = 8'hcc;
 buffer[1860] = 8'hcc;
 buffer[1861] = 8'h78;
 buffer[1862] = 8'h30;
 buffer[1863] = 8'hfc;
 buffer[1864] = 8'h38;
 buffer[1865] = 8'h6c;
 buffer[1866] = 8'hc6;
 buffer[1867] = 8'hfe;
 buffer[1868] = 8'hc6;
 buffer[1869] = 8'h6c;
 buffer[1870] = 8'h38;
 buffer[1871] = 8'h00;
 buffer[1872] = 8'h38;
 buffer[1873] = 8'h6c;
 buffer[1874] = 8'hc6;
 buffer[1875] = 8'hc6;
 buffer[1876] = 8'h6c;
 buffer[1877] = 8'h6c;
 buffer[1878] = 8'hee;
 buffer[1879] = 8'h00;
 buffer[1880] = 8'h1c;
 buffer[1881] = 8'h30;
 buffer[1882] = 8'h18;
 buffer[1883] = 8'h7c;
 buffer[1884] = 8'hcc;
 buffer[1885] = 8'hcc;
 buffer[1886] = 8'h78;
 buffer[1887] = 8'h00;
 buffer[1888] = 8'h00;
 buffer[1889] = 8'h00;
 buffer[1890] = 8'h7e;
 buffer[1891] = 8'hdb;
 buffer[1892] = 8'hdb;
 buffer[1893] = 8'h7e;
 buffer[1894] = 8'h00;
 buffer[1895] = 8'h00;
 buffer[1896] = 8'h06;
 buffer[1897] = 8'h0c;
 buffer[1898] = 8'h7e;
 buffer[1899] = 8'hdb;
 buffer[1900] = 8'hdb;
 buffer[1901] = 8'h7e;
 buffer[1902] = 8'h60;
 buffer[1903] = 8'hc0;
 buffer[1904] = 8'h38;
 buffer[1905] = 8'h60;
 buffer[1906] = 8'hc0;
 buffer[1907] = 8'hf8;
 buffer[1908] = 8'hc0;
 buffer[1909] = 8'h60;
 buffer[1910] = 8'h38;
 buffer[1911] = 8'h00;
 buffer[1912] = 8'h78;
 buffer[1913] = 8'hcc;
 buffer[1914] = 8'hcc;
 buffer[1915] = 8'hcc;
 buffer[1916] = 8'hcc;
 buffer[1917] = 8'hcc;
 buffer[1918] = 8'hcc;
 buffer[1919] = 8'h00;
 buffer[1920] = 8'h00;
 buffer[1921] = 8'hfc;
 buffer[1922] = 8'h00;
 buffer[1923] = 8'hfc;
 buffer[1924] = 8'h00;
 buffer[1925] = 8'hfc;
 buffer[1926] = 8'h00;
 buffer[1927] = 8'h00;
 buffer[1928] = 8'h30;
 buffer[1929] = 8'h30;
 buffer[1930] = 8'hfc;
 buffer[1931] = 8'h30;
 buffer[1932] = 8'h30;
 buffer[1933] = 8'h00;
 buffer[1934] = 8'hfc;
 buffer[1935] = 8'h00;
 buffer[1936] = 8'h60;
 buffer[1937] = 8'h30;
 buffer[1938] = 8'h18;
 buffer[1939] = 8'h30;
 buffer[1940] = 8'h60;
 buffer[1941] = 8'h00;
 buffer[1942] = 8'hfc;
 buffer[1943] = 8'h00;
 buffer[1944] = 8'h18;
 buffer[1945] = 8'h30;
 buffer[1946] = 8'h60;
 buffer[1947] = 8'h30;
 buffer[1948] = 8'h18;
 buffer[1949] = 8'h00;
 buffer[1950] = 8'hfc;
 buffer[1951] = 8'h00;
 buffer[1952] = 8'h0e;
 buffer[1953] = 8'h1b;
 buffer[1954] = 8'h1b;
 buffer[1955] = 8'h18;
 buffer[1956] = 8'h18;
 buffer[1957] = 8'h18;
 buffer[1958] = 8'h18;
 buffer[1959] = 8'h18;
 buffer[1960] = 8'h18;
 buffer[1961] = 8'h18;
 buffer[1962] = 8'h18;
 buffer[1963] = 8'h18;
 buffer[1964] = 8'h18;
 buffer[1965] = 8'hd8;
 buffer[1966] = 8'hd8;
 buffer[1967] = 8'h70;
 buffer[1968] = 8'h30;
 buffer[1969] = 8'h30;
 buffer[1970] = 8'h00;
 buffer[1971] = 8'hfc;
 buffer[1972] = 8'h00;
 buffer[1973] = 8'h30;
 buffer[1974] = 8'h30;
 buffer[1975] = 8'h00;
 buffer[1976] = 8'h00;
 buffer[1977] = 8'h76;
 buffer[1978] = 8'hdc;
 buffer[1979] = 8'h00;
 buffer[1980] = 8'h76;
 buffer[1981] = 8'hdc;
 buffer[1982] = 8'h00;
 buffer[1983] = 8'h00;
 buffer[1984] = 8'h38;
 buffer[1985] = 8'h6c;
 buffer[1986] = 8'h6c;
 buffer[1987] = 8'h38;
 buffer[1988] = 8'h00;
 buffer[1989] = 8'h00;
 buffer[1990] = 8'h00;
 buffer[1991] = 8'h00;
 buffer[1992] = 8'h00;
 buffer[1993] = 8'h00;
 buffer[1994] = 8'h00;
 buffer[1995] = 8'h18;
 buffer[1996] = 8'h18;
 buffer[1997] = 8'h00;
 buffer[1998] = 8'h00;
 buffer[1999] = 8'h00;
 buffer[2000] = 8'h00;
 buffer[2001] = 8'h00;
 buffer[2002] = 8'h00;
 buffer[2003] = 8'h00;
 buffer[2004] = 8'h18;
 buffer[2005] = 8'h00;
 buffer[2006] = 8'h00;
 buffer[2007] = 8'h00;
 buffer[2008] = 8'h0f;
 buffer[2009] = 8'h0c;
 buffer[2010] = 8'h0c;
 buffer[2011] = 8'h0c;
 buffer[2012] = 8'hec;
 buffer[2013] = 8'h6c;
 buffer[2014] = 8'h3c;
 buffer[2015] = 8'h1c;
 buffer[2016] = 8'h78;
 buffer[2017] = 8'h6c;
 buffer[2018] = 8'h6c;
 buffer[2019] = 8'h6c;
 buffer[2020] = 8'h6c;
 buffer[2021] = 8'h00;
 buffer[2022] = 8'h00;
 buffer[2023] = 8'h00;
 buffer[2024] = 8'h70;
 buffer[2025] = 8'h18;
 buffer[2026] = 8'h30;
 buffer[2027] = 8'h60;
 buffer[2028] = 8'h78;
 buffer[2029] = 8'h00;
 buffer[2030] = 8'h00;
 buffer[2031] = 8'h00;
 buffer[2032] = 8'h00;
 buffer[2033] = 8'h00;
 buffer[2034] = 8'h3c;
 buffer[2035] = 8'h3c;
 buffer[2036] = 8'h3c;
 buffer[2037] = 8'h3c;
 buffer[2038] = 8'h00;
 buffer[2039] = 8'h00;
 buffer[2040] = 8'h00;
 buffer[2041] = 8'h00;
 buffer[2042] = 8'h00;
 buffer[2043] = 8'h00;
 buffer[2044] = 8'h00;
 buffer[2045] = 8'h00;
 buffer[2046] = 8'h00;
 buffer[2047] = 8'h00;
end

endmodule

module M_gpu (
in_gpu_x,
in_gpu_y,
in_gpu_colour,
in_gpu_param0,
in_gpu_param1,
in_gpu_param2,
in_gpu_param3,
in_gpu_write,
in_blit1_writer_tile,
in_blit1_writer_line,
in_blit1_writer_bitmap,
in_vector_block_number,
in_vector_block_colour,
in_vector_block_xc,
in_vector_block_yc,
in_draw_vector,
in_vertices_writer_block,
in_vertices_writer_vertex,
in_vertices_writer_xdelta,
in_vertices_writer_ydelta,
in_vertices_writer_active,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_colour_write,
out_bitmap_write,
out_gpu_active,
out_vector_block_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_gpu_x;
input signed [10:0] in_gpu_y;
input  [7:0] in_gpu_colour;
input signed [10:0] in_gpu_param0;
input signed [10:0] in_gpu_param1;
input signed [10:0] in_gpu_param2;
input signed [10:0] in_gpu_param3;
input  [3:0] in_gpu_write;
input  [4:0] in_blit1_writer_tile;
input  [3:0] in_blit1_writer_line;
input  [15:0] in_blit1_writer_bitmap;
input  [4:0] in_vector_block_number;
input  [6:0] in_vector_block_colour;
input signed [10:0] in_vector_block_xc;
input signed [10:0] in_vector_block_yc;
input  [0:0] in_draw_vector;
input  [4:0] in_vertices_writer_block;
input  [5:0] in_vertices_writer_vertex;
input signed [5:0] in_vertices_writer_xdelta;
input signed [5:0] in_vertices_writer_ydelta;
input  [0:0] in_vertices_writer_active;
output signed [10:0] out_bitmap_x_write;
output signed [10:0] out_bitmap_y_write;
output  [6:0] out_bitmap_colour_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_gpu_active;
output  [0:0] out_vector_block_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [0:0] _w_vector_drawer_vector_block_active;
wire signed [10:0] _w_vector_drawer_gpu_x;
wire signed [10:0] _w_vector_drawer_gpu_y;
wire  [6:0] _w_vector_drawer_gpu_colour;
wire signed [10:0] _w_vector_drawer_gpu_param0;
wire signed [10:0] _w_vector_drawer_gpu_param1;
wire  [0:0] _w_vector_drawer_gpu_write;
wire _w_vector_drawer_done;
wire  [10:0] _w_GPUrectangle_bitmap_x_write;
wire  [10:0] _w_GPUrectangle_bitmap_y_write;
wire  [0:0] _w_GPUrectangle_bitmap_write;
wire  [0:0] _w_GPUrectangle_busy;
wire _w_GPUrectangle_done;
wire  [10:0] _w_GPUline_bitmap_x_write;
wire  [10:0] _w_GPUline_bitmap_y_write;
wire  [0:0] _w_GPUline_bitmap_write;
wire  [0:0] _w_GPUline_busy;
wire _w_GPUline_done;
wire  [10:0] _w_GPUcircle_bitmap_x_write;
wire  [10:0] _w_GPUcircle_bitmap_y_write;
wire  [0:0] _w_GPUcircle_bitmap_write;
wire  [0:0] _w_GPUcircle_busy;
wire _w_GPUcircle_done;
wire  [10:0] _w_GPUdisc_bitmap_x_write;
wire  [10:0] _w_GPUdisc_bitmap_y_write;
wire  [0:0] _w_GPUdisc_bitmap_write;
wire  [0:0] _w_GPUdisc_busy;
wire _w_GPUdisc_done;
wire  [10:0] _w_GPUtriangle_bitmap_x_write;
wire  [10:0] _w_GPUtriangle_bitmap_y_write;
wire  [0:0] _w_GPUtriangle_bitmap_write;
wire  [0:0] _w_GPUtriangle_busy;
wire _w_GPUtriangle_done;
wire  [10:0] _w_GPUblit_bitmap_x_write;
wire  [10:0] _w_GPUblit_bitmap_y_write;
wire  [0:0] _w_GPUblit_bitmap_write;
wire  [0:0] _w_GPUblit_busy;
wire  [8:0] _w_GPUblit_blit1tilemap_addr0;
wire _w_GPUblit_done;
wire  [10:0] _w_VECTORline_bitmap_x_write;
wire  [10:0] _w_VECTORline_bitmap_y_write;
wire  [0:0] _w_VECTORline_bitmap_write;
wire  [0:0] _w_VECTORline_busy;
wire _w_VECTORline_done;
wire  [15:0] _w_mem_blit1tilemap_rdata0;
wire  [7:0] _w_mem_characterGenerator8x8_rdata0;

reg  [0:0] _d_blit1tilemap_wenable1;
reg  [0:0] _q_blit1tilemap_wenable1;
reg  [15:0] _d_blit1tilemap_wdata1;
reg  [15:0] _q_blit1tilemap_wdata1;
reg  [8:0] _d_blit1tilemap_addr1;
reg  [8:0] _q_blit1tilemap_addr1;
reg  [10:0] _d_characterGenerator8x8_addr0;
reg  [10:0] _q_characterGenerator8x8_addr0;
reg  [0:0] _d_characterGenerator8x8_wenable1;
reg  [0:0] _q_characterGenerator8x8_wenable1;
reg  [7:0] _d_characterGenerator8x8_wdata1;
reg  [7:0] _q_characterGenerator8x8_wdata1;
reg  [10:0] _d_characterGenerator8x8_addr1;
reg  [10:0] _q_characterGenerator8x8_addr1;
reg  [6:0] _d_gpu_active_colour;
reg  [6:0] _q_gpu_active_colour;
reg signed [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg signed [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [6:0] _d_bitmap_colour_write,_q_bitmap_colour_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_gpu_active,_q_gpu_active;
reg  [0:0] _d_GPUrectangle_start,_q_GPUrectangle_start;
reg  [0:0] _d_GPUline_start,_q_GPUline_start;
reg  [0:0] _d_GPUcircle_start,_q_GPUcircle_start;
reg  [0:0] _d_GPUdisc_start,_q_GPUdisc_start;
reg  [0:0] _d_GPUtriangle_start,_q_GPUtriangle_start;
reg  [0:0] _d_GPUblit_start,_q_GPUblit_start;
reg  [0:0] _d_GPUblit_tilecharacter,_q_GPUblit_tilecharacter;
reg  [0:0] _d_VECTORline_start,_q_VECTORline_start;
reg  [4:0] _d_index,_q_index;
reg  _vector_drawer_run;
reg  _GPUrectangle_run;
reg  _GPUline_run;
reg  _GPUcircle_run;
reg  _GPUdisc_run;
reg  _GPUtriangle_run;
reg  _GPUblit_run;
reg  _VECTORline_run;
assign out_bitmap_x_write = _d_bitmap_x_write;
assign out_bitmap_y_write = _d_bitmap_y_write;
assign out_bitmap_colour_write = _d_bitmap_colour_write;
assign out_bitmap_write = _d_bitmap_write;
assign out_gpu_active = _q_gpu_active;
assign out_vector_block_active = _w_vector_drawer_vector_block_active;
assign out_done = (_q_index == 17);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_blit1tilemap_wenable1 <= 0;
_q_blit1tilemap_wdata1 <= 0;
_q_blit1tilemap_addr1 <= 0;
_q_characterGenerator8x8_addr0 <= 0;
_q_characterGenerator8x8_wenable1 <= 0;
_q_characterGenerator8x8_wdata1 <= 0;
_q_characterGenerator8x8_addr1 <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_blit1tilemap_wenable1 <= _d_blit1tilemap_wenable1;
_q_blit1tilemap_wdata1 <= _d_blit1tilemap_wdata1;
_q_blit1tilemap_addr1 <= _d_blit1tilemap_addr1;
_q_characterGenerator8x8_addr0 <= _d_characterGenerator8x8_addr0;
_q_characterGenerator8x8_wenable1 <= _d_characterGenerator8x8_wenable1;
_q_characterGenerator8x8_wdata1 <= _d_characterGenerator8x8_wdata1;
_q_characterGenerator8x8_addr1 <= _d_characterGenerator8x8_addr1;
_q_gpu_active_colour <= _d_gpu_active_colour;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_colour_write <= _d_bitmap_colour_write;
_q_bitmap_write <= _d_bitmap_write;
_q_gpu_active <= _d_gpu_active;
_q_index <= _d_index;
  end
_q_GPUrectangle_start <= _d_GPUrectangle_start;
_q_GPUline_start <= _d_GPUline_start;
_q_GPUcircle_start <= _d_GPUcircle_start;
_q_GPUdisc_start <= _d_GPUdisc_start;
_q_GPUtriangle_start <= _d_GPUtriangle_start;
_q_GPUblit_start <= _d_GPUblit_start;
_q_GPUblit_tilecharacter <= _d_GPUblit_tilecharacter;
_q_VECTORline_start <= _d_VECTORline_start;
end

M_vectors vector_drawer (
.in_vector_block_number(in_vector_block_number),
.in_vector_block_colour(in_vector_block_colour),
.in_vector_block_xc(in_vector_block_xc),
.in_vector_block_yc(in_vector_block_yc),
.in_draw_vector(in_draw_vector),
.in_vertices_writer_block(in_vertices_writer_block),
.in_vertices_writer_vertex(in_vertices_writer_vertex),
.in_vertices_writer_xdelta(in_vertices_writer_xdelta),
.in_vertices_writer_ydelta(in_vertices_writer_ydelta),
.in_vertices_writer_active(in_vertices_writer_active),
.in_gpu_active(_d_gpu_active),
.out_vector_block_active(_w_vector_drawer_vector_block_active),
.out_gpu_x(_w_vector_drawer_gpu_x),
.out_gpu_y(_w_vector_drawer_gpu_y),
.out_gpu_colour(_w_vector_drawer_gpu_colour),
.out_gpu_param0(_w_vector_drawer_gpu_param0),
.out_gpu_param1(_w_vector_drawer_gpu_param1),
.out_gpu_write(_w_vector_drawer_gpu_write),
.out_done(_w_vector_drawer_done),
.in_run(_vector_drawer_run),
.reset(reset),
.clock(clock)
);
M_rectangle GPUrectangle (
.in_x(in_gpu_x),
.in_y(in_gpu_y),
.in_param0(in_gpu_param0),
.in_param1(in_gpu_param1),
.in_start(_d_GPUrectangle_start),
.out_bitmap_x_write(_w_GPUrectangle_bitmap_x_write),
.out_bitmap_y_write(_w_GPUrectangle_bitmap_y_write),
.out_bitmap_write(_w_GPUrectangle_bitmap_write),
.out_busy(_w_GPUrectangle_busy),
.out_done(_w_GPUrectangle_done),
.in_run(_GPUrectangle_run),
.reset(reset),
.clock(clock)
);
M_line GPUline (
.in_x(in_gpu_x),
.in_y(in_gpu_y),
.in_param0(in_gpu_param0),
.in_param1(in_gpu_param1),
.in_start(_d_GPUline_start),
.out_bitmap_x_write(_w_GPUline_bitmap_x_write),
.out_bitmap_y_write(_w_GPUline_bitmap_y_write),
.out_bitmap_write(_w_GPUline_bitmap_write),
.out_busy(_w_GPUline_busy),
.out_done(_w_GPUline_done),
.in_run(_GPUline_run),
.reset(reset),
.clock(clock)
);
M_circle GPUcircle (
.in_x(in_gpu_x),
.in_y(in_gpu_y),
.in_param0(in_gpu_param0),
.in_start(_d_GPUcircle_start),
.out_bitmap_x_write(_w_GPUcircle_bitmap_x_write),
.out_bitmap_y_write(_w_GPUcircle_bitmap_y_write),
.out_bitmap_write(_w_GPUcircle_bitmap_write),
.out_busy(_w_GPUcircle_busy),
.out_done(_w_GPUcircle_done),
.in_run(_GPUcircle_run),
.reset(reset),
.clock(clock)
);
M_disc GPUdisc (
.in_x(in_gpu_x),
.in_y(in_gpu_y),
.in_param0(in_gpu_param0),
.in_start(_d_GPUdisc_start),
.out_bitmap_x_write(_w_GPUdisc_bitmap_x_write),
.out_bitmap_y_write(_w_GPUdisc_bitmap_y_write),
.out_bitmap_write(_w_GPUdisc_bitmap_write),
.out_busy(_w_GPUdisc_busy),
.out_done(_w_GPUdisc_done),
.in_run(_GPUdisc_run),
.reset(reset),
.clock(clock)
);
M_triangle GPUtriangle (
.in_x(in_gpu_x),
.in_y(in_gpu_y),
.in_param0(in_gpu_param0),
.in_param1(in_gpu_param1),
.in_param2(in_gpu_param2),
.in_param3(in_gpu_param3),
.in_start(_d_GPUtriangle_start),
.out_bitmap_x_write(_w_GPUtriangle_bitmap_x_write),
.out_bitmap_y_write(_w_GPUtriangle_bitmap_y_write),
.out_bitmap_write(_w_GPUtriangle_bitmap_write),
.out_busy(_w_GPUtriangle_busy),
.out_done(_w_GPUtriangle_done),
.in_run(_GPUtriangle_run),
.reset(reset),
.clock(clock)
);
M_blit #(
.BLIT1TILEMAP_ADDR0_WIDTH(9),
.BLIT1TILEMAP_ADDR0_INIT(0),
.BLIT1TILEMAP_ADDR0_SIGNED(0),
.BLIT1TILEMAP_RDATA0_WIDTH(16),
.BLIT1TILEMAP_RDATA0_INIT(0),
.BLIT1TILEMAP_RDATA0_SIGNED(0)
) GPUblit (
.in_x(in_gpu_x),
.in_y(in_gpu_y),
.in_param0(in_gpu_param0),
.in_param1(in_gpu_param1),
.in_start(_d_GPUblit_start),
.in_tilecharacter(_d_GPUblit_tilecharacter),
.in_blit1tilemap_rdata0(_w_mem_blit1tilemap_rdata0),
.out_bitmap_x_write(_w_GPUblit_bitmap_x_write),
.out_bitmap_y_write(_w_GPUblit_bitmap_y_write),
.out_bitmap_write(_w_GPUblit_bitmap_write),
.out_busy(_w_GPUblit_busy),
.out_blit1tilemap_addr0(_w_GPUblit_blit1tilemap_addr0),
.out_done(_w_GPUblit_done),
.in_run(_GPUblit_run),
.reset(reset),
.clock(clock)
);
M_line VECTORline (
.in_x(_w_vector_drawer_gpu_x),
.in_y(_w_vector_drawer_gpu_y),
.in_param0(_w_vector_drawer_gpu_param0),
.in_param1(_w_vector_drawer_gpu_param1),
.in_start(_d_VECTORline_start),
.out_bitmap_x_write(_w_VECTORline_bitmap_x_write),
.out_bitmap_y_write(_w_VECTORline_bitmap_y_write),
.out_bitmap_write(_w_VECTORline_bitmap_write),
.out_busy(_w_VECTORline_busy),
.out_done(_w_VECTORline_done),
.in_run(_VECTORline_run),
.reset(reset),
.clock(clock)
);

M_gpu_mem_blit1tilemap __mem__blit1tilemap(
.clock0(clock),
.clock1(clock),
.in_blit1tilemap_addr0(_w_GPUblit_blit1tilemap_addr0),
.in_blit1tilemap_wenable1(_d_blit1tilemap_wenable1),
.in_blit1tilemap_wdata1(_d_blit1tilemap_wdata1),
.in_blit1tilemap_addr1(_d_blit1tilemap_addr1),
.out_blit1tilemap_rdata0(_w_mem_blit1tilemap_rdata0)
);
M_gpu_mem_characterGenerator8x8 __mem__characterGenerator8x8(
.clock0(clock),
.clock1(clock),
.in_characterGenerator8x8_addr0(_d_characterGenerator8x8_addr0),
.in_characterGenerator8x8_wenable1(_d_characterGenerator8x8_wenable1),
.in_characterGenerator8x8_wdata1(_d_characterGenerator8x8_wdata1),
.in_characterGenerator8x8_addr1(_d_characterGenerator8x8_addr1),
.out_characterGenerator8x8_rdata0(_w_mem_characterGenerator8x8_rdata0)
);


always @* begin
_d_blit1tilemap_wenable1 = _q_blit1tilemap_wenable1;
_d_blit1tilemap_wdata1 = _q_blit1tilemap_wdata1;
_d_blit1tilemap_addr1 = _q_blit1tilemap_addr1;
_d_characterGenerator8x8_addr0 = _q_characterGenerator8x8_addr0;
_d_characterGenerator8x8_wenable1 = _q_characterGenerator8x8_wenable1;
_d_characterGenerator8x8_wdata1 = _q_characterGenerator8x8_wdata1;
_d_characterGenerator8x8_addr1 = _q_characterGenerator8x8_addr1;
_d_gpu_active_colour = _q_gpu_active_colour;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_colour_write = _q_bitmap_colour_write;
_d_bitmap_write = _q_bitmap_write;
_d_gpu_active = _q_gpu_active;
_d_GPUrectangle_start = _q_GPUrectangle_start;
_d_GPUline_start = _q_GPUline_start;
_d_GPUcircle_start = _q_GPUcircle_start;
_d_GPUdisc_start = _q_GPUdisc_start;
_d_GPUtriangle_start = _q_GPUtriangle_start;
_d_GPUblit_start = _q_GPUblit_start;
_d_GPUblit_tilecharacter = _q_GPUblit_tilecharacter;
_d_VECTORline_start = _q_VECTORline_start;
_d_index = _q_index;
_vector_drawer_run = 1;
_GPUrectangle_run = 1;
_GPUline_run = 1;
_GPUcircle_run = 1;
_GPUdisc_run = 1;
_GPUtriangle_run = 1;
_GPUblit_run = 1;
_VECTORline_run = 1;
// _always_pre
_d_blit1tilemap_addr1 = in_blit1_writer_tile*16+in_blit1_writer_line;
_d_blit1tilemap_wdata1 = in_blit1_writer_bitmap;
_d_blit1tilemap_wenable1 = 1;
_d_bitmap_write = 0;
_d_bitmap_colour_write = _q_gpu_active_colour;
_d_GPUrectangle_start = 0;
_d_GPUline_start = 0;
_d_GPUcircle_start = 0;
_d_GPUdisc_start = 0;
_d_GPUtriangle_start = 0;
_d_GPUblit_start = 0;
_d_VECTORline_start = 0;
_d_index = 17;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_blit1tilemap_wenable1 = 0;
_d_blit1tilemap_wdata1 = 0;
_d_blit1tilemap_addr1 = 0;
_d_characterGenerator8x8_addr0 = 0;
_d_characterGenerator8x8_wenable1 = 0;
_d_characterGenerator8x8_wdata1 = 0;
_d_characterGenerator8x8_addr1 = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (_w_vector_drawer_gpu_write) begin
// __block_5
// __block_7
_d_gpu_active_colour = _w_vector_drawer_gpu_colour;
_d_gpu_active = 1;
_d_VECTORline_start = 1;
_d_index = 3;
end else begin
// __block_6
// __block_14
_d_gpu_active_colour = in_gpu_colour;
  case (in_gpu_write)
  1: begin
// __block_16_case
// __block_17
_d_bitmap_x_write = in_gpu_x;
_d_bitmap_y_write = in_gpu_y;
_d_bitmap_write = 1;
// __block_18
_d_index = 1;
  end
  2: begin
// __block_19_case
// __block_20
_d_gpu_active = 1;
_d_GPUrectangle_start = 1;
_d_index = 5;
  end
  3: begin
// __block_27_case
// __block_28
_d_gpu_active = 1;
_d_GPUline_start = 1;
_d_index = 6;
  end
  4: begin
// __block_35_case
// __block_36
_d_gpu_active = 1;
_d_GPUcircle_start = 1;
_d_index = 7;
  end
  5: begin
// __block_43_case
// __block_44
_d_gpu_active = 1;
_d_GPUblit_start = 1;
_d_index = 8;
  end
  6: begin
// __block_51_case
// __block_52
_d_gpu_active = 1;
_d_GPUdisc_start = 1;
_d_index = 9;
  end
  7: begin
// __block_59_case
// __block_60
_d_gpu_active = 1;
_d_GPUtriangle_start = 1;
_d_index = 10;
  end
  default: begin
// __block_67_case
// __block_68
_d_gpu_active = 0;
// __block_69
_d_index = 1;
  end
endcase
end
end else begin
_d_index = 2;
end
end
3: begin
// __while__block_8
if (_w_VECTORline_busy) begin
// __block_9
// __block_11
_d_bitmap_x_write = _w_VECTORline_bitmap_x_write;
_d_bitmap_y_write = _w_VECTORline_bitmap_y_write;
_d_bitmap_write = _w_VECTORline_bitmap_write;
// __block_12
_d_index = 3;
end else begin
_d_index = 4;
end
end
5: begin
// __while__block_21
if (_w_GPUrectangle_busy) begin
// __block_22
// __block_24
_d_bitmap_x_write = _w_GPUrectangle_bitmap_x_write;
_d_bitmap_y_write = _w_GPUrectangle_bitmap_y_write;
_d_bitmap_write = _w_GPUrectangle_bitmap_write;
// __block_25
_d_index = 5;
end else begin
_d_index = 11;
end
end
6: begin
// __while__block_29
if (_w_GPUline_busy) begin
// __block_30
// __block_32
_d_bitmap_x_write = _w_GPUline_bitmap_x_write;
_d_bitmap_y_write = _w_GPUline_bitmap_y_write;
_d_bitmap_write = _w_GPUline_bitmap_write;
// __block_33
_d_index = 6;
end else begin
_d_index = 12;
end
end
7: begin
// __while__block_37
if (_w_GPUcircle_busy) begin
// __block_38
// __block_40
_d_bitmap_x_write = _w_GPUcircle_bitmap_x_write;
_d_bitmap_y_write = _w_GPUcircle_bitmap_y_write;
_d_bitmap_write = _w_GPUcircle_bitmap_write;
// __block_41
_d_index = 7;
end else begin
_d_index = 13;
end
end
8: begin
// __while__block_45
if (_w_GPUblit_busy) begin
// __block_46
// __block_48
_d_bitmap_x_write = _w_GPUblit_bitmap_x_write;
_d_bitmap_y_write = _w_GPUblit_bitmap_y_write;
_d_bitmap_write = _w_GPUblit_bitmap_write;
// __block_49
_d_index = 8;
end else begin
_d_index = 14;
end
end
9: begin
// __while__block_53
if (_w_GPUdisc_busy) begin
// __block_54
// __block_56
_d_bitmap_x_write = _w_GPUdisc_bitmap_x_write;
_d_bitmap_y_write = _w_GPUdisc_bitmap_y_write;
_d_bitmap_write = _w_GPUdisc_bitmap_write;
// __block_57
_d_index = 9;
end else begin
_d_index = 15;
end
end
10: begin
// __while__block_61
if (_w_GPUtriangle_busy) begin
// __block_62
// __block_64
_d_bitmap_x_write = _w_GPUtriangle_bitmap_x_write;
_d_bitmap_y_write = _w_GPUtriangle_bitmap_y_write;
_d_bitmap_write = _w_GPUtriangle_bitmap_write;
// __block_65
_d_index = 10;
end else begin
_d_index = 16;
end
end
2: begin
// __block_3
_d_index = 17;
end
4: begin
// __block_10
_d_gpu_active = 0;
// __block_13
_d_index = 1;
end
11: begin
// __block_23
_d_gpu_active = 0;
// __block_26
_d_index = 1;
end
12: begin
// __block_31
_d_gpu_active = 0;
// __block_34
_d_index = 1;
end
13: begin
// __block_39
_d_gpu_active = 0;
// __block_42
_d_index = 1;
end
14: begin
// __block_47
_d_gpu_active = 0;
// __block_50
_d_index = 1;
end
15: begin
// __block_55
_d_gpu_active = 0;
// __block_58
_d_index = 1;
end
16: begin
// __block_63
_d_gpu_active = 0;
// __block_66
_d_index = 1;
end
17: begin // end of gpu
end
default: begin 
_d_index = 17;
 end
endcase
end
endmodule


module M_rectangle (
in_x,
in_y,
in_param0,
in_param1,
in_start,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_write,
out_busy,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_x;
input signed [10:0] in_y;
input signed [10:0] in_param0;
input signed [10:0] in_param1;
input  [0:0] in_start;
output  [10:0] out_bitmap_x_write;
output  [10:0] out_bitmap_y_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_busy;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_gpu_active_x;
reg signed [10:0] _q_gpu_active_x;
reg signed [10:0] _d_gpu_active_y;
reg signed [10:0] _q_gpu_active_y;
reg signed [10:0] _d_gpu_x1;
reg signed [10:0] _q_gpu_x1;
reg signed [10:0] _d_gpu_max_x;
reg signed [10:0] _q_gpu_max_x;
reg signed [10:0] _d_gpu_max_y;
reg signed [10:0] _q_gpu_max_y;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg  [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_busy,_q_busy;
reg  [3:0] _d_index,_q_index;
assign out_bitmap_x_write = _d_bitmap_x_write;
assign out_bitmap_y_write = _d_bitmap_y_write;
assign out_bitmap_write = _d_bitmap_write;
assign out_busy = _q_busy;
assign out_done = (_q_index == 9);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_active <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_x1 <= _d_gpu_x1;
_q_gpu_max_x <= _d_gpu_max_x;
_q_gpu_max_y <= _d_gpu_max_y;
_q_active <= _d_active;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_write <= _d_bitmap_write;
_q_busy <= _d_busy;
_q_index <= _d_index;
  end
end




always @* begin
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_x1 = _q_gpu_x1;
_d_gpu_max_x = _q_gpu_max_x;
_d_gpu_max_y = _q_gpu_max_y;
_d_active = _q_active;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_write = _q_bitmap_write;
_d_busy = _q_busy;
_d_index = _q_index;
// _always_pre
_d_busy = in_start?1:_q_active;
_d_bitmap_write = 0;
_d_index = 9;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_active = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
_d_active = 1;
// __block_8_min
// __block_9
_d_gpu_active_x = (in_x<in_param0)?in_x:in_param0;
// __block_10
// __block_11
// __block_12_min
// __block_13
_d_gpu_active_y = (in_y<in_param1)?in_y:in_param1;
// __block_14
// __block_15
// __block_16_max
// __block_17
_d_gpu_max_x = (in_x>in_param0)?in_x:in_param0;
// __block_18
// __block_19
// __block_20_max
// __block_21
_d_gpu_max_y = (in_y>in_param1)?in_y:in_param1;
// __block_22
// __block_23
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_24
// __block_25_cropleft
// __block_26
_d_gpu_active_x = (_q_gpu_active_x<0)?0:_q_gpu_active_x;
// __block_27
// __block_28
// __block_29_cropleft
// __block_30
_d_gpu_x1 = (_d_gpu_active_x<0)?0:_d_gpu_active_x;
// __block_31
// __block_32
// __block_33_croptop
// __block_34
_d_gpu_active_y = (_q_gpu_active_y<0)?0:_q_gpu_active_y;
// __block_35
// __block_36
// __block_37_cropright
// __block_38
_d_gpu_max_x = (_q_gpu_max_x>639)?639:_q_gpu_max_x;
// __block_39
// __block_40
// __block_41_cropbottom
// __block_42
_d_gpu_max_y = (_q_gpu_max_y>479)?479:_q_gpu_max_y;
// __block_43
// __block_44
_d_index = 4;
end
2: begin
// __block_3
_d_index = 9;
end
4: begin
// __block_45
_d_index = 5;
end
5: begin
// __while__block_46
if (_q_gpu_active_y<=_q_gpu_max_y) begin
// __block_47
// __block_49
_d_bitmap_y_write = _q_gpu_active_y;
_d_index = 7;
end else begin
_d_index = 6;
end
end
7: begin
// __while__block_50
if (_q_gpu_active_x<=_q_gpu_max_x) begin
// __block_51
// __block_53
_d_bitmap_x_write = _q_gpu_active_x;
_d_bitmap_write = 1;
_d_gpu_active_x = _q_gpu_active_x+1;
// __block_54
_d_index = 7;
end else begin
_d_index = 8;
end
end
6: begin
// __block_48
_d_active = 0;
// __block_56
_d_index = 1;
end
8: begin
// __block_52
_d_gpu_active_x = _q_gpu_x1;
_d_gpu_active_y = _q_gpu_active_y+1;
// __block_55
_d_index = 5;
end
9: begin // end of rectangle
end
default: begin 
_d_index = 9;
 end
endcase
end
endmodule


module M_line (
in_x,
in_y,
in_param0,
in_param1,
in_start,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_write,
out_busy,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_x;
input signed [10:0] in_y;
input signed [10:0] in_param0;
input signed [10:0] in_param1;
input  [0:0] in_start;
output  [10:0] out_bitmap_x_write;
output  [10:0] out_bitmap_y_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_busy;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_gpu_active_x;
reg signed [10:0] _q_gpu_active_x;
reg signed [10:0] _d_gpu_active_y;
reg signed [10:0] _q_gpu_active_y;
reg signed [10:0] _d_gpu_dx;
reg signed [10:0] _q_gpu_dx;
reg signed [10:0] _d_gpu_dy;
reg signed [10:0] _q_gpu_dy;
reg signed [10:0] _d_gpu_sy;
reg signed [10:0] _q_gpu_sy;
reg signed [10:0] _d_gpu_numerator;
reg signed [10:0] _q_gpu_numerator;
reg signed [10:0] _d_gpu_numerator2;
reg signed [10:0] _q_gpu_numerator2;
reg signed [10:0] _d_gpu_count;
reg signed [10:0] _q_gpu_count;
reg signed [10:0] _d_gpu_max_count;
reg signed [10:0] _q_gpu_max_count;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg  [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_busy,_q_busy;
reg  [3:0] _d_index,_q_index;
assign out_bitmap_x_write = _d_bitmap_x_write;
assign out_bitmap_y_write = _d_bitmap_y_write;
assign out_bitmap_write = _d_bitmap_write;
assign out_busy = _q_busy;
assign out_done = (_q_index == 9);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_active <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_dx <= _d_gpu_dx;
_q_gpu_dy <= _d_gpu_dy;
_q_gpu_sy <= _d_gpu_sy;
_q_gpu_numerator <= _d_gpu_numerator;
_q_gpu_numerator2 <= _d_gpu_numerator2;
_q_gpu_count <= _d_gpu_count;
_q_gpu_max_count <= _d_gpu_max_count;
_q_active <= _d_active;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_write <= _d_bitmap_write;
_q_busy <= _d_busy;
_q_index <= _d_index;
  end
end




always @* begin
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_dx = _q_gpu_dx;
_d_gpu_dy = _q_gpu_dy;
_d_gpu_sy = _q_gpu_sy;
_d_gpu_numerator = _q_gpu_numerator;
_d_gpu_numerator2 = _q_gpu_numerator2;
_d_gpu_count = _q_gpu_count;
_d_gpu_max_count = _q_gpu_max_count;
_d_active = _q_active;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_write = _q_bitmap_write;
_d_busy = _q_busy;
_d_index = _q_index;
// _always_pre
_d_busy = in_start?1:_q_active;
_d_bitmap_write = 0;
_d_index = 9;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_active = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
_d_active = 1;
// __block_8_min
// __block_9
_d_gpu_active_x = (in_x<in_param0)?in_x:in_param0;
// __block_10
// __block_11
_d_gpu_active_y = (in_x<in_param0)?in_y:in_param1;
_d_gpu_sy = (in_x<in_param0)?((in_y<in_param1)?1:-1):((in_y<in_param1)?-1:1);
// __block_12_absdelta
// __block_13
_d_gpu_dx = (in_x<in_param0)?in_param0-in_x:in_x-in_param0;
// __block_14
// __block_15
// __block_16_absdelta
// __block_17
_d_gpu_dy = (in_y<in_param1)?in_param1-in_y:in_y-in_param1;
// __block_18
// __block_19
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_20
_d_gpu_count = 0;
_d_gpu_numerator = (_q_gpu_dx>_q_gpu_dy)?(_q_gpu_dx>>1):-(_q_gpu_dy>>1);
// __block_21_max
// __block_22
_d_gpu_max_count = (_q_gpu_dx>_q_gpu_dy)?_q_gpu_dx:_q_gpu_dy;
// __block_23
// __block_24
_d_index = 4;
end
2: begin
// __block_3
_d_index = 9;
end
4: begin
// __block_25
_d_index = 5;
end
5: begin
// __while__block_26
if (_q_gpu_count<=_q_gpu_max_count) begin
// __block_27
// __block_29
_d_bitmap_x_write = _q_gpu_active_x;
_d_bitmap_y_write = _q_gpu_active_y;
_d_bitmap_write = 1;
_d_gpu_numerator2 = _q_gpu_numerator;
_d_index = 7;
end else begin
_d_index = 6;
end
end
7: begin
// __block_30
if (_q_gpu_numerator2>(-_q_gpu_dx)) begin
// __block_31
// __block_33
_d_gpu_numerator = _q_gpu_numerator-_q_gpu_dy;
_d_gpu_active_x = _q_gpu_active_x+1;
// __block_34
end else begin
// __block_32
end
// __block_35
_d_index = 8;
end
6: begin
// __block_28
_d_active = 0;
// __block_43
_d_index = 1;
end
8: begin
// __block_36
if (_q_gpu_numerator2<_q_gpu_dy) begin
// __block_37
// __block_39
_d_gpu_numerator = _q_gpu_numerator+_q_gpu_dx;
_d_gpu_active_y = _q_gpu_active_y+_q_gpu_sy;
// __block_40
end else begin
// __block_38
end
// __block_41
_d_gpu_count = _q_gpu_count+1;
// __block_42
_d_index = 5;
end
9: begin // end of line
end
default: begin 
_d_index = 9;
 end
endcase
end
endmodule


module M_circle (
in_x,
in_y,
in_param0,
in_start,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_write,
out_busy,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_x;
input signed [10:0] in_y;
input signed [10:0] in_param0;
input  [0:0] in_start;
output  [10:0] out_bitmap_x_write;
output  [10:0] out_bitmap_y_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_busy;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_gpu_active_x;
reg signed [10:0] _q_gpu_active_x;
reg signed [10:0] _d_gpu_active_y;
reg signed [10:0] _q_gpu_active_y;
reg signed [10:0] _d_gpu_xc;
reg signed [10:0] _q_gpu_xc;
reg signed [10:0] _d_gpu_yc;
reg signed [10:0] _q_gpu_yc;
reg signed [10:0] _d_gpu_numerator;
reg signed [10:0] _q_gpu_numerator;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg  [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_busy,_q_busy;
reg  [3:0] _d_index,_q_index;
assign out_bitmap_x_write = _q_bitmap_x_write;
assign out_bitmap_y_write = _q_bitmap_y_write;
assign out_bitmap_write = _q_bitmap_write;
assign out_busy = _q_busy;
assign out_done = (_q_index == 14);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_active <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_xc <= _d_gpu_xc;
_q_gpu_yc <= _d_gpu_yc;
_q_gpu_numerator <= _d_gpu_numerator;
_q_active <= _d_active;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_write <= _d_bitmap_write;
_q_busy <= _d_busy;
_q_index <= _d_index;
  end
end




always @* begin
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_xc = _q_gpu_xc;
_d_gpu_yc = _q_gpu_yc;
_d_gpu_numerator = _q_gpu_numerator;
_d_active = _q_active;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_write = _q_bitmap_write;
_d_busy = _q_busy;
_d_index = _q_index;
// _always_pre
_d_busy = in_start?1:_q_active;
_d_bitmap_write = 0;
_d_index = 14;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_active = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
_d_active = 1;
_d_gpu_active_x = 0;
// __block_8_abs
// __block_9
_d_gpu_active_y = (in_param0<0)?-in_param0:in_param0;
// __block_10
// __block_11
// __block_12_copycoordinates
// __block_13
_d_gpu_xc = in_x;
_d_gpu_yc = in_y;
// __block_14
// __block_15
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_16
_d_gpu_numerator = 3-(2*_q_gpu_active_y);
_d_index = 4;
end
2: begin
// __block_3
_d_index = 14;
end
4: begin
// __block_17
_d_index = 5;
end
5: begin
// __while__block_18
if (_q_gpu_active_y>=_q_gpu_active_x) begin
// __block_19
// __block_21
_d_bitmap_x_write = _q_gpu_xc+_q_gpu_active_x;
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_active_y;
_d_bitmap_write = 1;
_d_index = 7;
end else begin
_d_index = 6;
end
end
7: begin
// __block_22
_d_bitmap_y_write = _q_gpu_yc-_q_gpu_active_y;
_d_bitmap_write = 1;
_d_index = 8;
end
6: begin
// __block_20
_d_active = 0;
// __block_37
_d_index = 1;
end
8: begin
// __block_23
_d_bitmap_x_write = _q_gpu_xc-_q_gpu_active_x;
_d_bitmap_write = 1;
_d_index = 9;
end
9: begin
// __block_24
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_active_y;
_d_bitmap_write = 1;
_d_index = 10;
end
10: begin
// __block_25
_d_bitmap_x_write = _q_gpu_xc+_q_gpu_active_y;
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_active_x;
_d_bitmap_write = 1;
_d_index = 11;
end
11: begin
// __block_26
_d_bitmap_y_write = _q_gpu_yc-_q_gpu_active_x;
_d_bitmap_write = 1;
_d_index = 12;
end
12: begin
// __block_27
_d_bitmap_x_write = _q_gpu_xc-_q_gpu_active_y;
_d_bitmap_write = 1;
_d_index = 13;
end
13: begin
// __block_28
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_active_x;
_d_bitmap_write = 1;
_d_gpu_active_x = _q_gpu_active_x+1;
if (_q_gpu_numerator>0) begin
// __block_29
// __block_31
_d_gpu_numerator = _q_gpu_numerator+4*(_d_gpu_active_x-_q_gpu_active_y)+10;
_d_gpu_active_y = _q_gpu_active_y-1;
// __block_32
end else begin
// __block_30
// __block_33
_d_gpu_numerator = _q_gpu_numerator+4*_d_gpu_active_x+6;
// __block_34
end
// __block_35
// __block_36
_d_index = 5;
end
14: begin // end of circle
end
default: begin 
_d_index = 14;
 end
endcase
end
endmodule


module M_disc (
in_x,
in_y,
in_param0,
in_start,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_write,
out_busy,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_x;
input signed [10:0] in_y;
input signed [10:0] in_param0;
input  [0:0] in_start;
output  [10:0] out_bitmap_x_write;
output  [10:0] out_bitmap_y_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_busy;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_gpu_active_x;
reg signed [10:0] _q_gpu_active_x;
reg signed [10:0] _d_gpu_active_y;
reg signed [10:0] _q_gpu_active_y;
reg signed [10:0] _d_gpu_xc;
reg signed [10:0] _q_gpu_xc;
reg signed [10:0] _d_gpu_yc;
reg signed [10:0] _q_gpu_yc;
reg signed [10:0] _d_gpu_numerator;
reg signed [10:0] _q_gpu_numerator;
reg signed [10:0] _d_gpu_count;
reg signed [10:0] _q_gpu_count;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg  [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_busy,_q_busy;
reg  [4:0] _d_index,_q_index;
assign out_bitmap_x_write = _q_bitmap_x_write;
assign out_bitmap_y_write = _q_bitmap_y_write;
assign out_bitmap_write = _q_bitmap_write;
assign out_busy = _q_busy;
assign out_done = (_q_index == 17);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_active <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_xc <= _d_gpu_xc;
_q_gpu_yc <= _d_gpu_yc;
_q_gpu_numerator <= _d_gpu_numerator;
_q_gpu_count <= _d_gpu_count;
_q_active <= _d_active;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_write <= _d_bitmap_write;
_q_busy <= _d_busy;
_q_index <= _d_index;
  end
end




always @* begin
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_xc = _q_gpu_xc;
_d_gpu_yc = _q_gpu_yc;
_d_gpu_numerator = _q_gpu_numerator;
_d_gpu_count = _q_gpu_count;
_d_active = _q_active;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_write = _q_bitmap_write;
_d_busy = _q_busy;
_d_index = _q_index;
// _always_pre
_d_busy = in_start?1:_q_active;
_d_bitmap_write = 0;
_d_index = 17;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_active = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
_d_active = 1;
_d_gpu_active_x = 0;
// __block_8_abs
// __block_9
_d_gpu_active_y = (in_param0<0)?-in_param0:in_param0;
// __block_10
// __block_11
// __block_12_copycoordinates
// __block_13
_d_gpu_xc = in_x;
_d_gpu_yc = in_y;
// __block_14
// __block_15
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_16
_d_gpu_active_y = (_q_gpu_active_y<4)?4:_q_gpu_active_y;
_d_index = 4;
end
2: begin
// __block_3
_d_index = 17;
end
4: begin
// __block_17
_d_gpu_count = _q_gpu_active_y;
_d_gpu_numerator = 3-(2*_q_gpu_active_y);
_d_index = 5;
end
5: begin
// __block_18
_d_index = 6;
end
6: begin
// __while__block_19
if (_q_gpu_active_y>=_q_gpu_active_x) begin
// __block_20
// __block_22
_d_index = 8;
end else begin
_d_index = 7;
end
end
8: begin
// __while__block_23
if (_q_gpu_count!=0) begin
// __block_24
// __block_26
_d_bitmap_x_write = _q_gpu_xc+_q_gpu_active_x;
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_count;
_d_bitmap_write = 1;
_d_index = 10;
end else begin
_d_index = 9;
end
end
7: begin
// __block_21
_d_bitmap_x_write = _q_gpu_xc;
_d_bitmap_y_write = _q_gpu_yc;
_d_bitmap_write = 1;
_d_active = 0;
// __block_43
_d_index = 1;
end
10: begin
// __block_27
_d_bitmap_y_write = _q_gpu_yc-_q_gpu_count;
_d_bitmap_write = 1;
_d_index = 11;
end
9: begin
// __block_25
_d_gpu_active_x = _q_gpu_active_x+1;
if (_q_gpu_numerator>0) begin
// __block_35
// __block_37
_d_gpu_numerator = _q_gpu_numerator+4*(_d_gpu_active_x-_q_gpu_active_y)+10;
_d_gpu_active_y = _q_gpu_active_y-1;
_d_gpu_count = _d_gpu_active_y-1;
// __block_38
end else begin
// __block_36
// __block_39
_d_gpu_numerator = _q_gpu_numerator+4*_d_gpu_active_x+6;
_d_gpu_count = _q_gpu_active_y;
// __block_40
end
// __block_41
// __block_42
_d_index = 6;
end
11: begin
// __block_28
_d_bitmap_x_write = _q_gpu_xc-_q_gpu_active_x;
_d_bitmap_write = 1;
_d_index = 12;
end
12: begin
// __block_29
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_count;
_d_bitmap_write = 1;
_d_index = 13;
end
13: begin
// __block_30
_d_bitmap_x_write = _q_gpu_xc+_q_gpu_count;
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_active_x;
_d_bitmap_write = 1;
_d_index = 14;
end
14: begin
// __block_31
_d_bitmap_y_write = _q_gpu_yc-_q_gpu_active_x;
_d_bitmap_write = 1;
_d_index = 15;
end
15: begin
// __block_32
_d_bitmap_x_write = _q_gpu_xc-_q_gpu_count;
_d_bitmap_write = 1;
_d_index = 16;
end
16: begin
// __block_33
_d_bitmap_y_write = _q_gpu_yc+_q_gpu_active_x;
_d_bitmap_write = 1;
_d_gpu_count = _q_gpu_count-1;
// __block_34
_d_index = 8;
end
17: begin // end of disc
end
default: begin 
_d_index = 17;
 end
endcase
end
endmodule


module M_triangle (
in_x,
in_y,
in_param0,
in_param1,
in_param2,
in_param3,
in_start,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_write,
out_busy,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_x;
input signed [10:0] in_y;
input signed [10:0] in_param0;
input signed [10:0] in_param1;
input signed [10:0] in_param2;
input signed [10:0] in_param3;
input  [0:0] in_start;
output  [10:0] out_bitmap_x_write;
output  [10:0] out_bitmap_y_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_busy;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_gpu_active_x;
reg signed [10:0] _q_gpu_active_x;
reg signed [10:0] _d_gpu_active_y;
reg signed [10:0] _q_gpu_active_y;
reg signed [10:0] _d_gpu_x1;
reg signed [10:0] _q_gpu_x1;
reg signed [10:0] _d_gpu_y1;
reg signed [10:0] _q_gpu_y1;
reg signed [10:0] _d_gpu_x2;
reg signed [10:0] _q_gpu_x2;
reg signed [10:0] _d_gpu_y2;
reg signed [10:0] _q_gpu_y2;
reg signed [10:0] _d_gpu_dx;
reg signed [10:0] _q_gpu_dx;
reg signed [10:0] _d_gpu_sx;
reg signed [10:0] _q_gpu_sx;
reg signed [10:0] _d_gpu_sy;
reg signed [10:0] _q_gpu_sy;
reg signed [10:0] _d_gpu_min_x;
reg signed [10:0] _q_gpu_min_x;
reg signed [10:0] _d_gpu_max_x;
reg signed [10:0] _q_gpu_max_x;
reg signed [10:0] _d_gpu_min_y;
reg signed [10:0] _q_gpu_min_y;
reg signed [10:0] _d_gpu_max_y;
reg signed [10:0] _q_gpu_max_y;
reg  [0:0] _d_gpu_count;
reg  [0:0] _q_gpu_count;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [0:0] _d_w0;
reg  [0:0] _q_w0;
reg  [0:0] _d_w1;
reg  [0:0] _q_w1;
reg  [0:0] _d_w2;
reg  [0:0] _q_w2;
reg  [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg  [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_busy,_q_busy;
reg  [3:0] _d_index,_q_index;
assign out_bitmap_x_write = _q_bitmap_x_write;
assign out_bitmap_y_write = _q_bitmap_y_write;
assign out_bitmap_write = _q_bitmap_write;
assign out_busy = _q_busy;
assign out_done = (_q_index == 14);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_active <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_x1 <= _d_gpu_x1;
_q_gpu_y1 <= _d_gpu_y1;
_q_gpu_x2 <= _d_gpu_x2;
_q_gpu_y2 <= _d_gpu_y2;
_q_gpu_dx <= _d_gpu_dx;
_q_gpu_sx <= _d_gpu_sx;
_q_gpu_sy <= _d_gpu_sy;
_q_gpu_min_x <= _d_gpu_min_x;
_q_gpu_max_x <= _d_gpu_max_x;
_q_gpu_min_y <= _d_gpu_min_y;
_q_gpu_max_y <= _d_gpu_max_y;
_q_gpu_count <= _d_gpu_count;
_q_active <= _d_active;
_q_w0 <= _d_w0;
_q_w1 <= _d_w1;
_q_w2 <= _d_w2;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_write <= _d_bitmap_write;
_q_busy <= _d_busy;
_q_index <= _d_index;
  end
end




always @* begin
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_x1 = _q_gpu_x1;
_d_gpu_y1 = _q_gpu_y1;
_d_gpu_x2 = _q_gpu_x2;
_d_gpu_y2 = _q_gpu_y2;
_d_gpu_dx = _q_gpu_dx;
_d_gpu_sx = _q_gpu_sx;
_d_gpu_sy = _q_gpu_sy;
_d_gpu_min_x = _q_gpu_min_x;
_d_gpu_max_x = _q_gpu_max_x;
_d_gpu_min_y = _q_gpu_min_y;
_d_gpu_max_y = _q_gpu_max_y;
_d_gpu_count = _q_gpu_count;
_d_active = _q_active;
_d_w0 = _q_w0;
_d_w1 = _q_w1;
_d_w2 = _q_w2;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_write = _q_bitmap_write;
_d_busy = _q_busy;
_d_index = _q_index;
// _always_pre
_d_busy = in_start?1:_q_active;
_d_bitmap_write = 0;
_d_index = 14;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_active = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
_d_active = 1;
// __block_8_copycoordinates
// __block_9
_d_gpu_active_x = in_x;
_d_gpu_active_y = in_y;
// __block_10
// __block_11
// __block_12_copycoordinates
// __block_13
_d_gpu_x1 = in_param0;
_d_gpu_y1 = in_param1;
// __block_14
// __block_15
// __block_16_copycoordinates
// __block_17
_d_gpu_x2 = in_param2;
_d_gpu_y2 = in_param3;
// __block_18
// __block_19
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_20
// __block_21_min3
// __block_22
_d_gpu_min_x = (_q_gpu_active_x<_q_gpu_x1)?(_q_gpu_active_x<_q_gpu_x2?_q_gpu_active_x:_q_gpu_x2):(_q_gpu_x1<_q_gpu_x2?_q_gpu_x1:_q_gpu_x2);
// __block_23
// __block_24
// __block_25_min3
// __block_26
_d_gpu_min_y = (_q_gpu_active_y<_q_gpu_y1)?(_q_gpu_active_y<_q_gpu_y2?_q_gpu_active_y:_q_gpu_y2):(_q_gpu_y1<_q_gpu_y2?_q_gpu_y1:_q_gpu_y2);
// __block_27
// __block_28
// __block_29_max3
// __block_30
_d_gpu_max_x = (_q_gpu_active_x>_q_gpu_x1)?(_q_gpu_active_x>_q_gpu_x2?_q_gpu_active_x:_q_gpu_x2):(_q_gpu_x1>_q_gpu_x2?_q_gpu_x1:_q_gpu_x2);
// __block_31
// __block_32
// __block_33_max3
// __block_34
_d_gpu_max_y = (_q_gpu_active_y>_q_gpu_y1)?(_q_gpu_active_y>_q_gpu_y2?_q_gpu_active_y:_q_gpu_y2):(_q_gpu_y1>_q_gpu_y2?_q_gpu_y1:_q_gpu_y2);
// __block_35
// __block_36
_d_index = 4;
end
2: begin
// __block_3
_d_index = 14;
end
4: begin
// __block_37
// __block_38_cropleft
// __block_39
_d_gpu_min_x = (_q_gpu_min_x<0)?0:_q_gpu_min_x;
// __block_40
// __block_41
// __block_42_cropright
// __block_43
_d_gpu_max_x = (_q_gpu_max_x>639)?639:_q_gpu_max_x;
// __block_44
// __block_45
// __block_46_croptop
// __block_47
_d_gpu_min_y = (_q_gpu_min_y<0)?0:_q_gpu_min_y;
// __block_48
// __block_49
// __block_50_cropbottom
// __block_51
_d_gpu_max_y = (_q_gpu_max_y>479)?479:_q_gpu_max_y;
// __block_52
// __block_53
_d_index = 5;
end
5: begin
// __block_54
if (_q_gpu_y1<_q_gpu_active_y) begin
// __block_55
// __block_57
// __block_58_swapcoordinates
// __block_59
_d_gpu_active_x = _q_gpu_x1;
_d_gpu_active_y = _q_gpu_y1;
_d_gpu_x1 = _d_gpu_active_x;
_d_gpu_y1 = _d_gpu_active_y;
// __block_60
// __block_61
// __block_62
end else begin
// __block_56
end
// __block_63
_d_index = 6;
end
6: begin
// __block_64
if (_q_gpu_y2<_q_gpu_active_y) begin
// __block_65
// __block_67
// __block_68_swapcoordinates
// __block_69
_d_gpu_active_x = _q_gpu_x2;
_d_gpu_active_y = _q_gpu_y2;
_d_gpu_x2 = _d_gpu_active_x;
_d_gpu_y2 = _d_gpu_active_y;
// __block_70
// __block_71
// __block_72
end else begin
// __block_66
end
// __block_73
_d_index = 7;
end
7: begin
// __block_74
if (_q_gpu_x1<_q_gpu_x2) begin
// __block_75
// __block_77
// __block_78_swapcoordinates
// __block_79
_d_gpu_x1 = _q_gpu_x2;
_d_gpu_y1 = _q_gpu_y2;
_d_gpu_x2 = _d_gpu_x1;
_d_gpu_y2 = _d_gpu_y1;
// __block_80
// __block_81
// __block_82
end else begin
// __block_76
end
// __block_83
_d_index = 8;
end
8: begin
// __block_84
// __block_85_copycoordinates
// __block_86
_d_gpu_sx = _q_gpu_min_x;
_d_gpu_sy = _q_gpu_min_y;
// __block_87
// __block_88
_d_gpu_dx = 1;
_d_gpu_count = 0;
_d_index = 9;
end
9: begin
// __block_89
_d_index = 10;
end
10: begin
// __while__block_90
if (_q_gpu_sy<=_q_gpu_max_y) begin
// __block_91
// __block_93
_d_w0 = ((_q_gpu_x2-_q_gpu_x1)*(_q_gpu_sy-_q_gpu_y1)-(_q_gpu_y2-_q_gpu_y1)*(_q_gpu_sx-_q_gpu_x1))>=0;
_d_w1 = ((_q_gpu_active_x-_q_gpu_x2)*(_q_gpu_sy-_q_gpu_y2)-(_q_gpu_active_y-_q_gpu_y2)*(_q_gpu_sx-_q_gpu_x2))>=0;
_d_w2 = ((_q_gpu_x1-_q_gpu_active_x)*(_q_gpu_sy-_q_gpu_active_y)-(_q_gpu_y1-_q_gpu_active_y)*(_q_gpu_sx-_q_gpu_active_x))>=0;
_d_index = 12;
end else begin
_d_index = 11;
end
end
12: begin
// __block_94
_d_bitmap_x_write = _q_gpu_sx;
_d_bitmap_y_write = _q_gpu_sy;
_d_bitmap_write = (_q_w0&&_q_w1&&_q_w2);
_d_gpu_count = (_q_w0&&_q_w1&&_q_w2)?1:_q_gpu_count;
_d_index = 13;
end
11: begin
// __block_92
_d_active = 0;
// __block_132
_d_index = 1;
end
13: begin
// __block_95
if (_q_gpu_count&&~(_q_w0&&_q_w1&&_q_w2)) begin
// __block_96
// __block_98
_d_gpu_count = 0;
_d_gpu_sy = _q_gpu_sy+1;
if ((_q_gpu_max_x-_q_gpu_sx)<(_q_gpu_sx-_q_gpu_min_x)) begin
// __block_99
// __block_101
_d_gpu_sx = _q_gpu_max_x;
_d_gpu_dx = -1;
// __block_102
end else begin
// __block_100
// __block_103
_d_gpu_sx = _q_gpu_min_x;
_d_gpu_dx = 1;
// __block_104
end
// __block_105
// __block_106
end else begin
// __block_97
// __block_107
  case (_q_gpu_dx)
  1: begin
// __block_109_case
// __block_110
if (_q_gpu_sx<_q_gpu_max_x) begin
// __block_111
// __block_113
_d_gpu_sx = _q_gpu_sx+1;
// __block_114
end else begin
// __block_112
// __block_115
_d_gpu_dx = -1;
_d_gpu_count = 0;
_d_gpu_sy = _q_gpu_sy+1;
// __block_116
end
// __block_117
// __block_118
  end
  default: begin
// __block_119_case
// __block_120
if (_q_gpu_sx>_q_gpu_min_x) begin
// __block_121
// __block_123
_d_gpu_sx = _q_gpu_sx-1;
// __block_124
end else begin
// __block_122
// __block_125
_d_gpu_dx = 1;
_d_gpu_count = 0;
_d_gpu_sy = _q_gpu_sy+1;
// __block_126
end
// __block_127
// __block_128
  end
endcase
// __block_108
// __block_129
end
// __block_130
// __block_131
_d_index = 10;
end
14: begin // end of triangle
end
default: begin 
_d_index = 14;
 end
endcase
end
endmodule


module M_blit #(
parameter BLIT1TILEMAP_ADDR0_WIDTH=1,parameter BLIT1TILEMAP_ADDR0_SIGNED=0,parameter BLIT1TILEMAP_ADDR0_INIT=0,
parameter BLIT1TILEMAP_RDATA0_WIDTH=1,parameter BLIT1TILEMAP_RDATA0_SIGNED=0,parameter BLIT1TILEMAP_RDATA0_INIT=0
) (
in_x,
in_y,
in_param0,
in_param1,
in_start,
in_tilecharacter,
in_blit1tilemap_rdata0,
out_bitmap_x_write,
out_bitmap_y_write,
out_bitmap_write,
out_busy,
out_blit1tilemap_addr0,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [10:0] in_x;
input signed [10:0] in_y;
input signed [10:0] in_param0;
input  [1:0] in_param1;
input  [0:0] in_start;
input  [0:0] in_tilecharacter;
input  [BLIT1TILEMAP_RDATA0_WIDTH-1:0] in_blit1tilemap_rdata0;
output  [10:0] out_bitmap_x_write;
output  [10:0] out_bitmap_y_write;
output  [0:0] out_bitmap_write;
output  [0:0] out_busy;
output  [BLIT1TILEMAP_ADDR0_WIDTH-1:0] out_blit1tilemap_addr0;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_gpu_active_x;
reg signed [10:0] _q_gpu_active_x;
reg signed [10:0] _d_gpu_active_y;
reg signed [10:0] _q_gpu_active_y;
reg signed [10:0] _d_gpu_x1;
reg signed [10:0] _q_gpu_x1;
reg signed [10:0] _d_gpu_y1;
reg signed [10:0] _q_gpu_y1;
reg signed [10:0] _d_gpu_max_x;
reg signed [10:0] _q_gpu_max_x;
reg signed [10:0] _d_gpu_max_y;
reg signed [10:0] _q_gpu_max_y;
reg  [7:0] _d_gpu_tile;
reg  [7:0] _q_gpu_tile;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [10:0] _d_bitmap_x_write,_q_bitmap_x_write;
reg  [10:0] _d_bitmap_y_write,_q_bitmap_y_write;
reg  [0:0] _d_bitmap_write,_q_bitmap_write;
reg  [0:0] _d_busy,_q_busy;
reg  [BLIT1TILEMAP_ADDR0_WIDTH-1:0] _d_blit1tilemap_addr0,_q_blit1tilemap_addr0;
reg  [3:0] _d_index,_q_index;
assign out_bitmap_x_write = _q_bitmap_x_write;
assign out_bitmap_y_write = _q_bitmap_y_write;
assign out_bitmap_write = _q_bitmap_write;
assign out_busy = _q_busy;
assign out_blit1tilemap_addr0 = _d_blit1tilemap_addr0;
assign out_done = (_q_index == 8);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_active <= 0;
_q_blit1tilemap_addr0 <= BLIT1TILEMAP_ADDR0_INIT;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_x1 <= _d_gpu_x1;
_q_gpu_y1 <= _d_gpu_y1;
_q_gpu_max_x <= _d_gpu_max_x;
_q_gpu_max_y <= _d_gpu_max_y;
_q_gpu_tile <= _d_gpu_tile;
_q_active <= _d_active;
_q_bitmap_x_write <= _d_bitmap_x_write;
_q_bitmap_y_write <= _d_bitmap_y_write;
_q_bitmap_write <= _d_bitmap_write;
_q_busy <= _d_busy;
_q_blit1tilemap_addr0 <= _d_blit1tilemap_addr0;
_q_index <= _d_index;
  end
end




always @* begin
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_x1 = _q_gpu_x1;
_d_gpu_y1 = _q_gpu_y1;
_d_gpu_max_x = _q_gpu_max_x;
_d_gpu_max_y = _q_gpu_max_y;
_d_gpu_tile = _q_gpu_tile;
_d_active = _q_active;
_d_bitmap_x_write = _q_bitmap_x_write;
_d_bitmap_y_write = _q_bitmap_y_write;
_d_bitmap_write = _q_bitmap_write;
_d_busy = _q_busy;
_d_blit1tilemap_addr0 = _q_blit1tilemap_addr0;
_d_index = _q_index;
// _always_pre
_d_blit1tilemap_addr0 = _q_gpu_tile*16+_q_gpu_active_y;
_d_busy = in_start?1:_q_active;
_d_bitmap_write = 0;
_d_index = 8;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_active = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
_d_active = 1;
_d_gpu_active_x = 0;
_d_gpu_active_y = 0;
// __block_8_copycoordinates
// __block_9
_d_gpu_x1 = in_x;
_d_gpu_y1 = in_y;
// __block_10
// __block_11
_d_gpu_max_x = 16;
_d_gpu_max_y = 16;
_d_gpu_tile = in_param0;
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_12
_d_index = 4;
end
2: begin
// __block_3
_d_index = 8;
end
4: begin
// __while__block_13
if (_q_gpu_active_y<_q_gpu_max_y) begin
// __block_14
// __block_16
_d_index = 6;
end else begin
_d_index = 5;
end
end
6: begin
// __while__block_17
if (_q_gpu_active_x<_q_gpu_max_x) begin
// __block_18
// __block_20
_d_bitmap_x_write = _q_gpu_x1+_q_gpu_active_x;
_d_bitmap_y_write = _q_gpu_y1+_q_gpu_active_y;
_d_bitmap_write = in_blit1tilemap_rdata0[15-_q_gpu_active_x+:1];
_d_gpu_active_x = _q_gpu_active_x+1;
// __block_21
_d_index = 6;
end else begin
_d_index = 7;
end
end
5: begin
// __block_15
_d_active = 0;
// __block_23
_d_index = 1;
end
7: begin
// __block_19
_d_gpu_active_x = 0;
_d_gpu_active_y = _q_gpu_active_y+1;
// __block_22
_d_index = 4;
end
8: begin // end of blit
end
default: begin 
_d_index = 8;
 end
endcase
end
endmodule


module M_vectors_mem_vertex(
input      [8:0]                in_vertex_addr0,
output reg  [12:0]     out_vertex_rdata0,
output reg  [12:0]     out_vertex_rdata1,
input      [0:0]             in_vertex_wenable1,
input      [12:0]                 in_vertex_wdata1,
input      [8:0]                in_vertex_addr1,
input      clock0,
input      clock1
);
reg  [12:0] buffer[511:0];
always @(posedge clock0) begin
  out_vertex_rdata0 <= buffer[in_vertex_addr0];
end
always @(posedge clock1) begin
  if (in_vertex_wenable1) begin
    buffer[in_vertex_addr1] <= in_vertex_wdata1;
  end
end

endmodule

module M_vectors (
in_vector_block_number,
in_vector_block_colour,
in_vector_block_xc,
in_vector_block_yc,
in_draw_vector,
in_vertices_writer_block,
in_vertices_writer_vertex,
in_vertices_writer_xdelta,
in_vertices_writer_ydelta,
in_vertices_writer_active,
in_gpu_active,
out_vector_block_active,
out_gpu_x,
out_gpu_y,
out_gpu_colour,
out_gpu_param0,
out_gpu_param1,
out_gpu_write,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [4:0] in_vector_block_number;
input  [6:0] in_vector_block_colour;
input signed [10:0] in_vector_block_xc;
input signed [10:0] in_vector_block_yc;
input  [0:0] in_draw_vector;
input  [4:0] in_vertices_writer_block;
input  [5:0] in_vertices_writer_vertex;
input signed [5:0] in_vertices_writer_xdelta;
input signed [5:0] in_vertices_writer_ydelta;
input  [0:0] in_vertices_writer_active;
input  [0:0] in_gpu_active;
output  [0:0] out_vector_block_active;
output signed [10:0] out_gpu_x;
output signed [10:0] out_gpu_y;
output  [6:0] out_gpu_colour;
output signed [10:0] out_gpu_param0;
output signed [10:0] out_gpu_param1;
output  [0:0] out_gpu_write;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [12:0] _w_mem_vertex_rdata0;
wire signed [10:0] _w_deltax;
wire signed [10:0] _w_deltay;

reg  [8:0] _d_vertex_addr0;
reg  [8:0] _q_vertex_addr0;
reg  [0:0] _d_vertex_wenable1;
reg  [0:0] _q_vertex_wenable1;
reg  [12:0] _d_vertex_wdata1;
reg  [12:0] _q_vertex_wdata1;
reg  [8:0] _d_vertex_addr1;
reg  [8:0] _q_vertex_addr1;
reg  [4:0] _d_block_number;
reg  [4:0] _q_block_number;
reg  [4:0] _d_vertices_number;
reg  [4:0] _q_vertices_number;
reg signed [10:0] _d_start_x;
reg signed [10:0] _q_start_x;
reg signed [10:0] _d_start_y;
reg signed [10:0] _q_start_y;
reg  [0:0] _d_vector_block_active,_q_vector_block_active;
reg signed [10:0] _d_gpu_x,_q_gpu_x;
reg signed [10:0] _d_gpu_y,_q_gpu_y;
reg  [6:0] _d_gpu_colour,_q_gpu_colour;
reg signed [10:0] _d_gpu_param0,_q_gpu_param0;
reg signed [10:0] _d_gpu_param1,_q_gpu_param1;
reg  [0:0] _d_gpu_write,_q_gpu_write;
reg  [3:0] _d_index,_q_index;
assign out_vector_block_active = _q_vector_block_active;
assign out_gpu_x = _q_gpu_x;
assign out_gpu_y = _q_gpu_y;
assign out_gpu_colour = _q_gpu_colour;
assign out_gpu_param0 = _q_gpu_param0;
assign out_gpu_param1 = _q_gpu_param1;
assign out_gpu_write = _q_gpu_write;
assign out_done = (_q_index == 10);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_vertex_addr0 <= 0;
_q_vertex_wenable1 <= 0;
_q_vertex_wdata1 <= 0;
_q_vertex_addr1 <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_vertex_addr0 <= _d_vertex_addr0;
_q_vertex_wenable1 <= _d_vertex_wenable1;
_q_vertex_wdata1 <= _d_vertex_wdata1;
_q_vertex_addr1 <= _d_vertex_addr1;
_q_block_number <= _d_block_number;
_q_vertices_number <= _d_vertices_number;
_q_start_x <= _d_start_x;
_q_start_y <= _d_start_y;
_q_vector_block_active <= _d_vector_block_active;
_q_gpu_x <= _d_gpu_x;
_q_gpu_y <= _d_gpu_y;
_q_gpu_colour <= _d_gpu_colour;
_q_gpu_param0 <= _d_gpu_param0;
_q_gpu_param1 <= _d_gpu_param1;
_q_gpu_write <= _d_gpu_write;
_q_index <= _d_index;
  end
end


M_vectors_mem_vertex __mem__vertex(
.clock0(clock),
.clock1(clock),
.in_vertex_addr0(_d_vertex_addr0),
.in_vertex_wenable1(_d_vertex_wenable1),
.in_vertex_wdata1(_d_vertex_wdata1),
.in_vertex_addr1(_d_vertex_addr1),
.out_vertex_rdata0(_w_mem_vertex_rdata0)
);

assign _w_deltay = {{6{_w_mem_vertex_rdata0[5+:1]}},_w_mem_vertex_rdata0[0+:5]};
assign _w_deltax = {{6{_w_mem_vertex_rdata0[11+:1]}},_w_mem_vertex_rdata0[6+:5]};

always @* begin
_d_vertex_addr0 = _q_vertex_addr0;
_d_vertex_wenable1 = _q_vertex_wenable1;
_d_vertex_wdata1 = _q_vertex_wdata1;
_d_vertex_addr1 = _q_vertex_addr1;
_d_block_number = _q_block_number;
_d_vertices_number = _q_vertices_number;
_d_start_x = _q_start_x;
_d_start_y = _q_start_y;
_d_vector_block_active = _q_vector_block_active;
_d_gpu_x = _q_gpu_x;
_d_gpu_y = _q_gpu_y;
_d_gpu_colour = _q_gpu_colour;
_d_gpu_param0 = _q_gpu_param0;
_d_gpu_param1 = _q_gpu_param1;
_d_gpu_write = _q_gpu_write;
_d_index = _q_index;
// _always_pre
_d_vertex_addr0 = _q_block_number*16+_q_vertices_number;
_d_vertex_addr1 = in_vertices_writer_block*16+in_vertices_writer_vertex;
_d_vertex_wdata1 = {in_vertices_writer_active,$unsigned(in_vertices_writer_xdelta),$unsigned(in_vertices_writer_ydelta)};
_d_vertex_wenable1 = 1;
_d_gpu_write = 0;
_d_index = 10;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_vertex_addr0 = 0;
_d_vertex_wenable1 = 0;
_d_vertex_wdata1 = 0;
_d_vertex_addr1 = 0;
// --
_d_vector_block_active = 0;
_d_vertices_number = 0;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_draw_vector) begin
// __block_5
// __block_7
_d_block_number = in_vector_block_number;
_d_gpu_colour = in_vector_block_colour;
_d_vertices_number = 0;
_d_vector_block_active = 1;
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_8
// __block_9_deltacoordinates
// __block_10
_d_start_x = in_vector_block_xc+_w_deltax;
_d_start_y = in_vector_block_yc+_w_deltay;
// __block_11
// __block_12
_d_vertices_number = 1;
_d_index = 4;
end
2: begin
// __block_3
_d_index = 10;
end
4: begin
// __block_13
_d_index = 5;
end
5: begin
// __while__block_14
if (_w_mem_vertex_rdata0[12+:1]&&(_q_vertices_number<16)) begin
// __block_15
// __block_17
// __block_18_copycoordinates
// __block_19
_d_gpu_x = _q_start_x;
_d_gpu_y = _q_start_y;
// __block_20
// __block_21
// __block_22_deltacoordinates
// __block_23
_d_gpu_param0 = in_vector_block_xc+_w_deltax;
_d_gpu_param1 = in_vector_block_yc+_w_deltay;
// __block_24
// __block_25
_d_index = 7;
end else begin
_d_index = 6;
end
end
7: begin
// __while__block_26
if (in_gpu_active) begin
// __block_27
// __block_29
// __block_30
_d_index = 7;
end else begin
_d_index = 8;
end
end
6: begin
// __block_16
_d_vector_block_active = 0;
// __block_37
_d_index = 1;
end
8: begin
// __block_28
_d_gpu_write = 1;
// __block_31_deltacoordinates
// __block_32
_d_start_x = in_vector_block_xc+_w_deltax;
_d_start_y = in_vector_block_yc+_w_deltay;
// __block_33
// __block_34
_d_vertices_number = _q_vertices_number+1;
_d_index = 9;
end
9: begin
// __block_35
// __block_36
_d_index = 5;
end
10: begin // end of vectors
end
default: begin 
_d_index = 10;
 end
endcase
end
endmodule


module M_background (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_staticGenerator,
in_backgroundcolour,
in_backgroundcolour_alt,
in_backgroundcolour_mode,
in_background_write,
out_pix_red,
out_pix_green,
out_pix_blue,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [15:0] in_staticGenerator;
input  [5:0] in_backgroundcolour;
input  [5:0] in_backgroundcolour_alt;
input  [3:0] in_backgroundcolour_mode;
input  [2:0] in_background_write;
output  [1:0] out_pix_red;
output  [1:0] out_pix_green;
output  [1:0] out_pix_blue;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
reg signed [9:0] _t_dotpos;
reg signed [1:0] _t_speed;

reg  [5:0] _d_background;
reg  [5:0] _q_background;
reg  [5:0] _d_background_alt;
reg  [5:0] _q_background_alt;
reg  [3:0] _d_background_mode;
reg  [3:0] _q_background_mode;
reg signed [11:0] _d_rand_x;
reg signed [11:0] _q_rand_x;
reg signed [31:0] _d_frame;
reg signed [31:0] _q_frame;
reg  [1:0] _d_pix_red,_q_pix_red;
reg  [1:0] _d_pix_green,_q_pix_green;
reg  [1:0] _d_pix_blue,_q_pix_blue;
reg  [1:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_background <= 0;
_q_background_alt <= 0;
_q_background_mode <= 0;
_q_rand_x <= 0;
_q_frame <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_background <= _d_background;
_q_background_alt <= _d_background_alt;
_q_background_mode <= _d_background_mode;
_q_rand_x <= _d_rand_x;
_q_frame <= _d_frame;
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_index <= _d_index;
  end
end




always @* begin
_d_background = _q_background;
_d_background_alt = _q_background_alt;
_d_background_mode = _q_background_mode;
_d_rand_x = _q_rand_x;
_d_frame = _q_frame;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_index = _q_index;
_t_dotpos = 0;
_t_speed = 0;
// _always_pre
_d_pix_red = _q_background[4+:2];
_d_pix_green = _q_background[2+:2];
_d_pix_blue = _q_background[0+:2];
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_background = 0;
_d_background_alt = 0;
_d_background_mode = 0;
_t_dotpos = 0;
_t_speed = 0;
_d_rand_x = 0;
_d_frame = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (in_background_write)
  1: begin
// __block_6_case
// __block_7
_d_background = in_backgroundcolour;
// __block_8
  end
  2: begin
// __block_9_case
// __block_10
_d_background_alt = in_backgroundcolour_alt;
// __block_11
  end
  3: begin
// __block_12_case
// __block_13
_d_background_mode = in_backgroundcolour_mode;
// __block_14
  end
endcase
// __block_5
_d_frame = ((in_pix_x==639)&&(in_pix_y==470))?_q_frame+1:_q_frame;
if (in_pix_active) begin
// __block_15
// __block_17
  case (_d_background_mode)
  1: begin
// __block_19_case
// __block_20
  case ({in_pix_x[0+:1],in_pix_y[0+:1]})
  2'b00: begin
// __block_22_case
// __block_23
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_24
  end
  2'b01: begin
// __block_25_case
// __block_26
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_27
  end
  2'b10: begin
// __block_28_case
// __block_29
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_30
  end
  2'b11: begin
// __block_31_case
// __block_32
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_33
  end
endcase
// __block_21
// __block_34
  end
  2: begin
// __block_35_case
// __block_36
  case ({in_pix_x[1+:1],in_pix_y[1+:1]})
  2'b00: begin
// __block_38_case
// __block_39
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_40
  end
  2'b01: begin
// __block_41_case
// __block_42
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_43
  end
  2'b10: begin
// __block_44_case
// __block_45
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_46
  end
  2'b11: begin
// __block_47_case
// __block_48
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_49
  end
endcase
// __block_37
// __block_50
  end
  3: begin
// __block_51_case
// __block_52
  case ({in_pix_x[2+:1],in_pix_y[2+:1]})
  2'b00: begin
// __block_54_case
// __block_55
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_56
  end
  2'b01: begin
// __block_57_case
// __block_58
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_59
  end
  2'b10: begin
// __block_60_case
// __block_61
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_62
  end
  2'b11: begin
// __block_63_case
// __block_64
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_65
  end
endcase
// __block_53
// __block_66
  end
  4: begin
// __block_67_case
// __block_68
  case ({in_pix_x[3+:1],in_pix_y[3+:1]})
  2'b00: begin
// __block_70_case
// __block_71
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_72
  end
  2'b01: begin
// __block_73_case
// __block_74
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_75
  end
  2'b10: begin
// __block_76_case
// __block_77
_d_pix_red = _d_background_alt[4+:2];
_d_pix_green = _d_background_alt[2+:2];
_d_pix_blue = _d_background_alt[0+:2];
// __block_78
  end
  2'b11: begin
// __block_79_case
// __block_80
_d_pix_red = _d_background[4+:2];
_d_pix_green = _d_background[2+:2];
_d_pix_blue = _d_background[0+:2];
// __block_81
  end
endcase
// __block_69
// __block_82
  end
  5: begin
// __block_83_case
// __block_84
  case (in_pix_y[6+:3])
  3'b000: begin
// __block_86_case
// __block_87
_d_pix_red = 2;
// __block_88
  end
  3'b001: begin
// __block_89_case
// __block_90
_d_pix_red = 3;
// __block_91
  end
  3'b010: begin
// __block_92_case
// __block_93
_d_pix_red = 3;
_d_pix_green = 2;
// __block_94
  end
  3'b011: begin
// __block_95_case
// __block_96
_d_pix_red = 3;
_d_pix_green = 3;
// __block_97
  end
  3'b100: begin
// __block_98_case
// __block_99
_d_pix_green = 3;
// __block_100
  end
  3'b101: begin
// __block_101_case
// __block_102
_d_pix_blue = 3;
// __block_103
  end
  3'b110: begin
// __block_104_case
// __block_105
_d_pix_red = 1;
_d_pix_blue = 2;
// __block_106
  end
  3'b111: begin
// __block_107_case
// __block_108
_d_pix_red = 1;
_d_pix_green = 2;
_d_pix_blue = 3;
// __block_109
  end
endcase
// __block_85
// __block_110
  end
  6: begin
// __block_111_case
// __block_112
_d_pix_red = in_staticGenerator[0+:2];
_d_pix_green = in_staticGenerator[0+:2];
_d_pix_blue = in_staticGenerator[0+:2];
// __block_113
  end
  7: begin
// __block_114_case
// __block_115
_d_rand_x = (in_pix_x==0)?1:_q_rand_x*31421+6927;
_t_speed = _d_rand_x[10+:2];
_t_dotpos = (_d_frame>>_t_speed)+_d_rand_x;
_d_pix_red = (in_pix_y==_t_dotpos)?_d_background[4+:2]:_d_background_alt[4+:2];
_d_pix_green = (in_pix_y==_t_dotpos)?_d_background[2+:2]:_d_background_alt[2+:2];
_d_pix_blue = (in_pix_y==_t_dotpos)?_d_background[0+:2]:_d_background_alt[0+:2];
// __block_116
  end
endcase
// __block_18
// __block_117
end else begin
// __block_16
end
// __block_118
// __block_119
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of background
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_sprite_layer_mem_tiles_0(
input      [6:0]                in_tiles_0_addr0,
output reg  [15:0]     out_tiles_0_rdata0,
output reg  [15:0]     out_tiles_0_rdata1,
input      [0:0]             in_tiles_0_wenable1,
input      [15:0]                 in_tiles_0_wdata1,
input      [6:0]                in_tiles_0_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_0_rdata0 <= buffer[in_tiles_0_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_0_wenable1) begin
    buffer[in_tiles_0_addr1] <= in_tiles_0_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_1(
input      [6:0]                in_tiles_1_addr0,
output reg  [15:0]     out_tiles_1_rdata0,
output reg  [15:0]     out_tiles_1_rdata1,
input      [0:0]             in_tiles_1_wenable1,
input      [15:0]                 in_tiles_1_wdata1,
input      [6:0]                in_tiles_1_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_1_rdata0 <= buffer[in_tiles_1_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_1_wenable1) begin
    buffer[in_tiles_1_addr1] <= in_tiles_1_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_2(
input      [6:0]                in_tiles_2_addr0,
output reg  [15:0]     out_tiles_2_rdata0,
output reg  [15:0]     out_tiles_2_rdata1,
input      [0:0]             in_tiles_2_wenable1,
input      [15:0]                 in_tiles_2_wdata1,
input      [6:0]                in_tiles_2_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_2_rdata0 <= buffer[in_tiles_2_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_2_wenable1) begin
    buffer[in_tiles_2_addr1] <= in_tiles_2_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_3(
input      [6:0]                in_tiles_3_addr0,
output reg  [15:0]     out_tiles_3_rdata0,
output reg  [15:0]     out_tiles_3_rdata1,
input      [0:0]             in_tiles_3_wenable1,
input      [15:0]                 in_tiles_3_wdata1,
input      [6:0]                in_tiles_3_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_3_rdata0 <= buffer[in_tiles_3_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_3_wenable1) begin
    buffer[in_tiles_3_addr1] <= in_tiles_3_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_4(
input      [6:0]                in_tiles_4_addr0,
output reg  [15:0]     out_tiles_4_rdata0,
output reg  [15:0]     out_tiles_4_rdata1,
input      [0:0]             in_tiles_4_wenable1,
input      [15:0]                 in_tiles_4_wdata1,
input      [6:0]                in_tiles_4_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_4_rdata0 <= buffer[in_tiles_4_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_4_wenable1) begin
    buffer[in_tiles_4_addr1] <= in_tiles_4_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_5(
input      [6:0]                in_tiles_5_addr0,
output reg  [15:0]     out_tiles_5_rdata0,
output reg  [15:0]     out_tiles_5_rdata1,
input      [0:0]             in_tiles_5_wenable1,
input      [15:0]                 in_tiles_5_wdata1,
input      [6:0]                in_tiles_5_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_5_rdata0 <= buffer[in_tiles_5_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_5_wenable1) begin
    buffer[in_tiles_5_addr1] <= in_tiles_5_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_6(
input      [6:0]                in_tiles_6_addr0,
output reg  [15:0]     out_tiles_6_rdata0,
output reg  [15:0]     out_tiles_6_rdata1,
input      [0:0]             in_tiles_6_wenable1,
input      [15:0]                 in_tiles_6_wdata1,
input      [6:0]                in_tiles_6_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_6_rdata0 <= buffer[in_tiles_6_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_6_wenable1) begin
    buffer[in_tiles_6_addr1] <= in_tiles_6_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_7(
input      [6:0]                in_tiles_7_addr0,
output reg  [15:0]     out_tiles_7_rdata0,
output reg  [15:0]     out_tiles_7_rdata1,
input      [0:0]             in_tiles_7_wenable1,
input      [15:0]                 in_tiles_7_wdata1,
input      [6:0]                in_tiles_7_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_7_rdata0 <= buffer[in_tiles_7_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_7_wenable1) begin
    buffer[in_tiles_7_addr1] <= in_tiles_7_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_8(
input      [6:0]                in_tiles_8_addr0,
output reg  [15:0]     out_tiles_8_rdata0,
output reg  [15:0]     out_tiles_8_rdata1,
input      [0:0]             in_tiles_8_wenable1,
input      [15:0]                 in_tiles_8_wdata1,
input      [6:0]                in_tiles_8_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_8_rdata0 <= buffer[in_tiles_8_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_8_wenable1) begin
    buffer[in_tiles_8_addr1] <= in_tiles_8_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_9(
input      [6:0]                in_tiles_9_addr0,
output reg  [15:0]     out_tiles_9_rdata0,
output reg  [15:0]     out_tiles_9_rdata1,
input      [0:0]             in_tiles_9_wenable1,
input      [15:0]                 in_tiles_9_wdata1,
input      [6:0]                in_tiles_9_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_9_rdata0 <= buffer[in_tiles_9_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_9_wenable1) begin
    buffer[in_tiles_9_addr1] <= in_tiles_9_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_10(
input      [6:0]                in_tiles_10_addr0,
output reg  [15:0]     out_tiles_10_rdata0,
output reg  [15:0]     out_tiles_10_rdata1,
input      [0:0]             in_tiles_10_wenable1,
input      [15:0]                 in_tiles_10_wdata1,
input      [6:0]                in_tiles_10_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_10_rdata0 <= buffer[in_tiles_10_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_10_wenable1) begin
    buffer[in_tiles_10_addr1] <= in_tiles_10_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_11(
input      [6:0]                in_tiles_11_addr0,
output reg  [15:0]     out_tiles_11_rdata0,
output reg  [15:0]     out_tiles_11_rdata1,
input      [0:0]             in_tiles_11_wenable1,
input      [15:0]                 in_tiles_11_wdata1,
input      [6:0]                in_tiles_11_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_11_rdata0 <= buffer[in_tiles_11_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_11_wenable1) begin
    buffer[in_tiles_11_addr1] <= in_tiles_11_wdata1;
  end
end

endmodule

module M_sprite_layer_mem_tiles_12(
input      [6:0]                in_tiles_12_addr0,
output reg  [15:0]     out_tiles_12_rdata0,
output reg  [15:0]     out_tiles_12_rdata1,
input      [0:0]             in_tiles_12_wenable1,
input      [15:0]                 in_tiles_12_wdata1,
input      [6:0]                in_tiles_12_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[127:0];
always @(posedge clock0) begin
  out_tiles_12_rdata0 <= buffer[in_tiles_12_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_12_wenable1) begin
    buffer[in_tiles_12_addr1] <= in_tiles_12_wdata1;
  end
end

endmodule

module M_sprite_layer (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_sprite_set_number,
in_sprite_set_active,
in_sprite_set_double,
in_sprite_set_colour,
in_sprite_set_x,
in_sprite_set_y,
in_sprite_set_tile,
in_sprite_layer_write,
in_sprite_update,
in_collision_layer_1,
in_collision_layer_2,
in_collision_layer_3,
in_sprite_writer_sprite,
in_sprite_writer_line,
in_sprite_writer_bitmap,
in_sprite_writer_active,
out_pix_red,
out_pix_green,
out_pix_blue,
out_sprite_layer_display,
out_sprite_read_active,
out_sprite_read_double,
out_sprite_read_colour,
out_sprite_read_x,
out_sprite_read_y,
out_sprite_read_tile,
out_collision_0,
out_collision_1,
out_collision_2,
out_collision_3,
out_collision_4,
out_collision_5,
out_collision_6,
out_collision_7,
out_collision_8,
out_collision_9,
out_collision_10,
out_collision_11,
out_collision_12,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [3:0] in_sprite_set_number;
input  [0:0] in_sprite_set_active;
input  [0:0] in_sprite_set_double;
input  [5:0] in_sprite_set_colour;
input signed [10:0] in_sprite_set_x;
input signed [10:0] in_sprite_set_y;
input  [2:0] in_sprite_set_tile;
input  [3:0] in_sprite_layer_write;
input  [15:0] in_sprite_update;
input  [0:0] in_collision_layer_1;
input  [0:0] in_collision_layer_2;
input  [0:0] in_collision_layer_3;
input  [3:0] in_sprite_writer_sprite;
input  [6:0] in_sprite_writer_line;
input  [15:0] in_sprite_writer_bitmap;
input  [0:0] in_sprite_writer_active;
output  [1:0] out_pix_red;
output  [1:0] out_pix_green;
output  [1:0] out_pix_blue;
output  [0:0] out_sprite_layer_display;
output  [0:0] out_sprite_read_active;
output  [0:0] out_sprite_read_double;
output  [5:0] out_sprite_read_colour;
output signed [10:0] out_sprite_read_x;
output signed [10:0] out_sprite_read_y;
output  [2:0] out_sprite_read_tile;
output  [15:0] out_collision_0;
output  [15:0] out_collision_1;
output  [15:0] out_collision_2;
output  [15:0] out_collision_3;
output  [15:0] out_collision_4;
output  [15:0] out_collision_5;
output  [15:0] out_collision_6;
output  [15:0] out_collision_7;
output  [15:0] out_collision_8;
output  [15:0] out_collision_9;
output  [15:0] out_collision_10;
output  [15:0] out_collision_11;
output  [15:0] out_collision_12;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [15:0] _w_mem_tiles_0_rdata0;
wire  [15:0] _w_mem_tiles_1_rdata0;
wire  [15:0] _w_mem_tiles_2_rdata0;
wire  [15:0] _w_mem_tiles_3_rdata0;
wire  [15:0] _w_mem_tiles_4_rdata0;
wire  [15:0] _w_mem_tiles_5_rdata0;
wire  [15:0] _w_mem_tiles_6_rdata0;
wire  [15:0] _w_mem_tiles_7_rdata0;
wire  [15:0] _w_mem_tiles_8_rdata0;
wire  [15:0] _w_mem_tiles_9_rdata0;
wire  [15:0] _w_mem_tiles_10_rdata0;
wire  [15:0] _w_mem_tiles_11_rdata0;
wire  [15:0] _w_mem_tiles_12_rdata0;
reg  [6:0] _t_tiles_0_addr0;
reg  [0:0] _t_tiles_0_wenable1;
reg  [15:0] _t_tiles_0_wdata1;
reg  [6:0] _t_tiles_0_addr1;
reg  [6:0] _t_tiles_1_addr0;
reg  [0:0] _t_tiles_1_wenable1;
reg  [15:0] _t_tiles_1_wdata1;
reg  [6:0] _t_tiles_1_addr1;
reg  [6:0] _t_tiles_2_addr0;
reg  [0:0] _t_tiles_2_wenable1;
reg  [15:0] _t_tiles_2_wdata1;
reg  [6:0] _t_tiles_2_addr1;
reg  [6:0] _t_tiles_3_addr0;
reg  [0:0] _t_tiles_3_wenable1;
reg  [15:0] _t_tiles_3_wdata1;
reg  [6:0] _t_tiles_3_addr1;
reg  [6:0] _t_tiles_4_addr0;
reg  [0:0] _t_tiles_4_wenable1;
reg  [15:0] _t_tiles_4_wdata1;
reg  [6:0] _t_tiles_4_addr1;
reg  [6:0] _t_tiles_5_addr0;
reg  [0:0] _t_tiles_5_wenable1;
reg  [15:0] _t_tiles_5_wdata1;
reg  [6:0] _t_tiles_5_addr1;
reg  [6:0] _t_tiles_6_addr0;
reg  [0:0] _t_tiles_6_wenable1;
reg  [15:0] _t_tiles_6_wdata1;
reg  [6:0] _t_tiles_6_addr1;
reg  [6:0] _t_tiles_7_addr0;
reg  [0:0] _t_tiles_7_wenable1;
reg  [15:0] _t_tiles_7_wdata1;
reg  [6:0] _t_tiles_7_addr1;
reg  [6:0] _t_tiles_8_addr0;
reg  [0:0] _t_tiles_8_wenable1;
reg  [15:0] _t_tiles_8_wdata1;
reg  [6:0] _t_tiles_8_addr1;
reg  [6:0] _t_tiles_9_addr0;
reg  [0:0] _t_tiles_9_wenable1;
reg  [15:0] _t_tiles_9_wdata1;
reg  [6:0] _t_tiles_9_addr1;
reg  [6:0] _t_tiles_10_addr0;
reg  [0:0] _t_tiles_10_wenable1;
reg  [15:0] _t_tiles_10_wdata1;
reg  [6:0] _t_tiles_10_addr1;
reg  [6:0] _t_tiles_11_addr0;
reg  [0:0] _t_tiles_11_wenable1;
reg  [15:0] _t_tiles_11_wdata1;
reg  [6:0] _t_tiles_11_addr1;
reg  [6:0] _t_tiles_12_addr0;
reg  [0:0] _t_tiles_12_wenable1;
reg  [15:0] _t_tiles_12_wdata1;
reg  [6:0] _t_tiles_12_addr1;
wire  [5:0] _w_spritesize_0;
wire  [0:0] _w_xinrange_0;
wire  [0:0] _w_yinrange_0;
wire  [0:0] _w_pix_visible_0;
wire  [5:0] _w_spritesize_1;
wire  [0:0] _w_xinrange_1;
wire  [0:0] _w_yinrange_1;
wire  [0:0] _w_pix_visible_1;
wire  [5:0] _w_spritesize_2;
wire  [0:0] _w_xinrange_2;
wire  [0:0] _w_yinrange_2;
wire  [0:0] _w_pix_visible_2;
wire  [5:0] _w_spritesize_3;
wire  [0:0] _w_xinrange_3;
wire  [0:0] _w_yinrange_3;
wire  [0:0] _w_pix_visible_3;
wire  [5:0] _w_spritesize_4;
wire  [0:0] _w_xinrange_4;
wire  [0:0] _w_yinrange_4;
wire  [0:0] _w_pix_visible_4;
wire  [5:0] _w_spritesize_5;
wire  [0:0] _w_xinrange_5;
wire  [0:0] _w_yinrange_5;
wire  [0:0] _w_pix_visible_5;
wire  [5:0] _w_spritesize_6;
wire  [0:0] _w_xinrange_6;
wire  [0:0] _w_yinrange_6;
wire  [0:0] _w_pix_visible_6;
wire  [5:0] _w_spritesize_7;
wire  [0:0] _w_xinrange_7;
wire  [0:0] _w_yinrange_7;
wire  [0:0] _w_pix_visible_7;
wire  [5:0] _w_spritesize_8;
wire  [0:0] _w_xinrange_8;
wire  [0:0] _w_yinrange_8;
wire  [0:0] _w_pix_visible_8;
wire  [5:0] _w_spritesize_9;
wire  [0:0] _w_xinrange_9;
wire  [0:0] _w_yinrange_9;
wire  [0:0] _w_pix_visible_9;
wire  [5:0] _w_spritesize_10;
wire  [0:0] _w_xinrange_10;
wire  [0:0] _w_yinrange_10;
wire  [0:0] _w_pix_visible_10;
wire  [5:0] _w_spritesize_11;
wire  [0:0] _w_xinrange_11;
wire  [0:0] _w_yinrange_11;
wire  [0:0] _w_pix_visible_11;
wire  [5:0] _w_spritesize_12;
wire  [0:0] _w_xinrange_12;
wire  [0:0] _w_yinrange_12;
wire  [0:0] _w_pix_visible_12;
wire signed [10:0] _w_deltax;
wire signed [10:0] _w_deltay;
wire signed [10:0] _w_sprite_offscreen_negative;
wire signed [10:0] _w_sprite_to_negative;
wire  [0:0] _w_sprite_offscreen_x;
wire  [0:0] _w_sprite_offscreen_y;

reg  [0:0] _d_sprite_active[12:0];
reg  [0:0] _q_sprite_active[12:0];
reg  [0:0] _d_sprite_double[12:0];
reg  [0:0] _q_sprite_double[12:0];
reg signed [10:0] _d_sprite_x[12:0];
reg signed [10:0] _q_sprite_x[12:0];
reg signed [10:0] _d_sprite_y[12:0];
reg signed [10:0] _q_sprite_y[12:0];
reg  [5:0] _d_sprite_colour[12:0];
reg  [5:0] _q_sprite_colour[12:0];
reg  [2:0] _d_sprite_tile_number[12:0];
reg  [2:0] _q_sprite_tile_number[12:0];
reg  [0:0] _d_output_collisions;
reg  [0:0] _q_output_collisions;
reg  [15:0] _d_detect_collision_0;
reg  [15:0] _q_detect_collision_0;
reg  [15:0] _d_detect_collision_1;
reg  [15:0] _q_detect_collision_1;
reg  [15:0] _d_detect_collision_2;
reg  [15:0] _q_detect_collision_2;
reg  [15:0] _d_detect_collision_3;
reg  [15:0] _q_detect_collision_3;
reg  [15:0] _d_detect_collision_4;
reg  [15:0] _q_detect_collision_4;
reg  [15:0] _d_detect_collision_5;
reg  [15:0] _q_detect_collision_5;
reg  [15:0] _d_detect_collision_6;
reg  [15:0] _q_detect_collision_6;
reg  [15:0] _d_detect_collision_7;
reg  [15:0] _q_detect_collision_7;
reg  [15:0] _d_detect_collision_8;
reg  [15:0] _q_detect_collision_8;
reg  [15:0] _d_detect_collision_9;
reg  [15:0] _q_detect_collision_9;
reg  [15:0] _d_detect_collision_10;
reg  [15:0] _q_detect_collision_10;
reg  [15:0] _d_detect_collision_11;
reg  [15:0] _q_detect_collision_11;
reg  [15:0] _d_detect_collision_12;
reg  [15:0] _q_detect_collision_12;
reg  [1:0] _d_pix_red,_q_pix_red;
reg  [1:0] _d_pix_green,_q_pix_green;
reg  [1:0] _d_pix_blue,_q_pix_blue;
reg  [0:0] _d_sprite_layer_display,_q_sprite_layer_display;
reg  [0:0] _d_sprite_read_active,_q_sprite_read_active;
reg  [0:0] _d_sprite_read_double,_q_sprite_read_double;
reg  [5:0] _d_sprite_read_colour,_q_sprite_read_colour;
reg signed [10:0] _d_sprite_read_x,_q_sprite_read_x;
reg signed [10:0] _d_sprite_read_y,_q_sprite_read_y;
reg  [2:0] _d_sprite_read_tile,_q_sprite_read_tile;
reg  [15:0] _d_collision_0,_q_collision_0;
reg  [15:0] _d_collision_1,_q_collision_1;
reg  [15:0] _d_collision_2,_q_collision_2;
reg  [15:0] _d_collision_3,_q_collision_3;
reg  [15:0] _d_collision_4,_q_collision_4;
reg  [15:0] _d_collision_5,_q_collision_5;
reg  [15:0] _d_collision_6,_q_collision_6;
reg  [15:0] _d_collision_7,_q_collision_7;
reg  [15:0] _d_collision_8,_q_collision_8;
reg  [15:0] _d_collision_9,_q_collision_9;
reg  [15:0] _d_collision_10,_q_collision_10;
reg  [15:0] _d_collision_11,_q_collision_11;
reg  [15:0] _d_collision_12,_q_collision_12;
reg  [1:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_sprite_layer_display = _d_sprite_layer_display;
assign out_sprite_read_active = _q_sprite_read_active;
assign out_sprite_read_double = _q_sprite_read_double;
assign out_sprite_read_colour = _q_sprite_read_colour;
assign out_sprite_read_x = _q_sprite_read_x;
assign out_sprite_read_y = _q_sprite_read_y;
assign out_sprite_read_tile = _q_sprite_read_tile;
assign out_collision_0 = _q_collision_0;
assign out_collision_1 = _q_collision_1;
assign out_collision_2 = _q_collision_2;
assign out_collision_3 = _q_collision_3;
assign out_collision_4 = _q_collision_4;
assign out_collision_5 = _q_collision_5;
assign out_collision_6 = _q_collision_6;
assign out_collision_7 = _q_collision_7;
assign out_collision_8 = _q_collision_8;
assign out_collision_9 = _q_collision_9;
assign out_collision_10 = _q_collision_10;
assign out_collision_11 = _q_collision_11;
assign out_collision_12 = _q_collision_12;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_output_collisions <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_sprite_active[0] <= _d_sprite_active[0];
_q_sprite_active[1] <= _d_sprite_active[1];
_q_sprite_active[2] <= _d_sprite_active[2];
_q_sprite_active[3] <= _d_sprite_active[3];
_q_sprite_active[4] <= _d_sprite_active[4];
_q_sprite_active[5] <= _d_sprite_active[5];
_q_sprite_active[6] <= _d_sprite_active[6];
_q_sprite_active[7] <= _d_sprite_active[7];
_q_sprite_active[8] <= _d_sprite_active[8];
_q_sprite_active[9] <= _d_sprite_active[9];
_q_sprite_active[10] <= _d_sprite_active[10];
_q_sprite_active[11] <= _d_sprite_active[11];
_q_sprite_active[12] <= _d_sprite_active[12];
_q_sprite_double[0] <= _d_sprite_double[0];
_q_sprite_double[1] <= _d_sprite_double[1];
_q_sprite_double[2] <= _d_sprite_double[2];
_q_sprite_double[3] <= _d_sprite_double[3];
_q_sprite_double[4] <= _d_sprite_double[4];
_q_sprite_double[5] <= _d_sprite_double[5];
_q_sprite_double[6] <= _d_sprite_double[6];
_q_sprite_double[7] <= _d_sprite_double[7];
_q_sprite_double[8] <= _d_sprite_double[8];
_q_sprite_double[9] <= _d_sprite_double[9];
_q_sprite_double[10] <= _d_sprite_double[10];
_q_sprite_double[11] <= _d_sprite_double[11];
_q_sprite_double[12] <= _d_sprite_double[12];
_q_sprite_x[0] <= _d_sprite_x[0];
_q_sprite_x[1] <= _d_sprite_x[1];
_q_sprite_x[2] <= _d_sprite_x[2];
_q_sprite_x[3] <= _d_sprite_x[3];
_q_sprite_x[4] <= _d_sprite_x[4];
_q_sprite_x[5] <= _d_sprite_x[5];
_q_sprite_x[6] <= _d_sprite_x[6];
_q_sprite_x[7] <= _d_sprite_x[7];
_q_sprite_x[8] <= _d_sprite_x[8];
_q_sprite_x[9] <= _d_sprite_x[9];
_q_sprite_x[10] <= _d_sprite_x[10];
_q_sprite_x[11] <= _d_sprite_x[11];
_q_sprite_x[12] <= _d_sprite_x[12];
_q_sprite_y[0] <= _d_sprite_y[0];
_q_sprite_y[1] <= _d_sprite_y[1];
_q_sprite_y[2] <= _d_sprite_y[2];
_q_sprite_y[3] <= _d_sprite_y[3];
_q_sprite_y[4] <= _d_sprite_y[4];
_q_sprite_y[5] <= _d_sprite_y[5];
_q_sprite_y[6] <= _d_sprite_y[6];
_q_sprite_y[7] <= _d_sprite_y[7];
_q_sprite_y[8] <= _d_sprite_y[8];
_q_sprite_y[9] <= _d_sprite_y[9];
_q_sprite_y[10] <= _d_sprite_y[10];
_q_sprite_y[11] <= _d_sprite_y[11];
_q_sprite_y[12] <= _d_sprite_y[12];
_q_sprite_colour[0] <= _d_sprite_colour[0];
_q_sprite_colour[1] <= _d_sprite_colour[1];
_q_sprite_colour[2] <= _d_sprite_colour[2];
_q_sprite_colour[3] <= _d_sprite_colour[3];
_q_sprite_colour[4] <= _d_sprite_colour[4];
_q_sprite_colour[5] <= _d_sprite_colour[5];
_q_sprite_colour[6] <= _d_sprite_colour[6];
_q_sprite_colour[7] <= _d_sprite_colour[7];
_q_sprite_colour[8] <= _d_sprite_colour[8];
_q_sprite_colour[9] <= _d_sprite_colour[9];
_q_sprite_colour[10] <= _d_sprite_colour[10];
_q_sprite_colour[11] <= _d_sprite_colour[11];
_q_sprite_colour[12] <= _d_sprite_colour[12];
_q_sprite_tile_number[0] <= _d_sprite_tile_number[0];
_q_sprite_tile_number[1] <= _d_sprite_tile_number[1];
_q_sprite_tile_number[2] <= _d_sprite_tile_number[2];
_q_sprite_tile_number[3] <= _d_sprite_tile_number[3];
_q_sprite_tile_number[4] <= _d_sprite_tile_number[4];
_q_sprite_tile_number[5] <= _d_sprite_tile_number[5];
_q_sprite_tile_number[6] <= _d_sprite_tile_number[6];
_q_sprite_tile_number[7] <= _d_sprite_tile_number[7];
_q_sprite_tile_number[8] <= _d_sprite_tile_number[8];
_q_sprite_tile_number[9] <= _d_sprite_tile_number[9];
_q_sprite_tile_number[10] <= _d_sprite_tile_number[10];
_q_sprite_tile_number[11] <= _d_sprite_tile_number[11];
_q_sprite_tile_number[12] <= _d_sprite_tile_number[12];
_q_output_collisions <= _d_output_collisions;
_q_detect_collision_0 <= _d_detect_collision_0;
_q_detect_collision_1 <= _d_detect_collision_1;
_q_detect_collision_2 <= _d_detect_collision_2;
_q_detect_collision_3 <= _d_detect_collision_3;
_q_detect_collision_4 <= _d_detect_collision_4;
_q_detect_collision_5 <= _d_detect_collision_5;
_q_detect_collision_6 <= _d_detect_collision_6;
_q_detect_collision_7 <= _d_detect_collision_7;
_q_detect_collision_8 <= _d_detect_collision_8;
_q_detect_collision_9 <= _d_detect_collision_9;
_q_detect_collision_10 <= _d_detect_collision_10;
_q_detect_collision_11 <= _d_detect_collision_11;
_q_detect_collision_12 <= _d_detect_collision_12;
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_sprite_layer_display <= _d_sprite_layer_display;
_q_sprite_read_active <= _d_sprite_read_active;
_q_sprite_read_double <= _d_sprite_read_double;
_q_sprite_read_colour <= _d_sprite_read_colour;
_q_sprite_read_x <= _d_sprite_read_x;
_q_sprite_read_y <= _d_sprite_read_y;
_q_sprite_read_tile <= _d_sprite_read_tile;
_q_collision_0 <= _d_collision_0;
_q_collision_1 <= _d_collision_1;
_q_collision_2 <= _d_collision_2;
_q_collision_3 <= _d_collision_3;
_q_collision_4 <= _d_collision_4;
_q_collision_5 <= _d_collision_5;
_q_collision_6 <= _d_collision_6;
_q_collision_7 <= _d_collision_7;
_q_collision_8 <= _d_collision_8;
_q_collision_9 <= _d_collision_9;
_q_collision_10 <= _d_collision_10;
_q_collision_11 <= _d_collision_11;
_q_collision_12 <= _d_collision_12;
_q_index <= _d_index;
  end
end


M_sprite_layer_mem_tiles_0 __mem__tiles_0(
.clock0(clock),
.clock1(clock),
.in_tiles_0_addr0(_t_tiles_0_addr0),
.in_tiles_0_wenable1(_t_tiles_0_wenable1),
.in_tiles_0_wdata1(_t_tiles_0_wdata1),
.in_tiles_0_addr1(_t_tiles_0_addr1),
.out_tiles_0_rdata0(_w_mem_tiles_0_rdata0)
);
M_sprite_layer_mem_tiles_1 __mem__tiles_1(
.clock0(clock),
.clock1(clock),
.in_tiles_1_addr0(_t_tiles_1_addr0),
.in_tiles_1_wenable1(_t_tiles_1_wenable1),
.in_tiles_1_wdata1(_t_tiles_1_wdata1),
.in_tiles_1_addr1(_t_tiles_1_addr1),
.out_tiles_1_rdata0(_w_mem_tiles_1_rdata0)
);
M_sprite_layer_mem_tiles_2 __mem__tiles_2(
.clock0(clock),
.clock1(clock),
.in_tiles_2_addr0(_t_tiles_2_addr0),
.in_tiles_2_wenable1(_t_tiles_2_wenable1),
.in_tiles_2_wdata1(_t_tiles_2_wdata1),
.in_tiles_2_addr1(_t_tiles_2_addr1),
.out_tiles_2_rdata0(_w_mem_tiles_2_rdata0)
);
M_sprite_layer_mem_tiles_3 __mem__tiles_3(
.clock0(clock),
.clock1(clock),
.in_tiles_3_addr0(_t_tiles_3_addr0),
.in_tiles_3_wenable1(_t_tiles_3_wenable1),
.in_tiles_3_wdata1(_t_tiles_3_wdata1),
.in_tiles_3_addr1(_t_tiles_3_addr1),
.out_tiles_3_rdata0(_w_mem_tiles_3_rdata0)
);
M_sprite_layer_mem_tiles_4 __mem__tiles_4(
.clock0(clock),
.clock1(clock),
.in_tiles_4_addr0(_t_tiles_4_addr0),
.in_tiles_4_wenable1(_t_tiles_4_wenable1),
.in_tiles_4_wdata1(_t_tiles_4_wdata1),
.in_tiles_4_addr1(_t_tiles_4_addr1),
.out_tiles_4_rdata0(_w_mem_tiles_4_rdata0)
);
M_sprite_layer_mem_tiles_5 __mem__tiles_5(
.clock0(clock),
.clock1(clock),
.in_tiles_5_addr0(_t_tiles_5_addr0),
.in_tiles_5_wenable1(_t_tiles_5_wenable1),
.in_tiles_5_wdata1(_t_tiles_5_wdata1),
.in_tiles_5_addr1(_t_tiles_5_addr1),
.out_tiles_5_rdata0(_w_mem_tiles_5_rdata0)
);
M_sprite_layer_mem_tiles_6 __mem__tiles_6(
.clock0(clock),
.clock1(clock),
.in_tiles_6_addr0(_t_tiles_6_addr0),
.in_tiles_6_wenable1(_t_tiles_6_wenable1),
.in_tiles_6_wdata1(_t_tiles_6_wdata1),
.in_tiles_6_addr1(_t_tiles_6_addr1),
.out_tiles_6_rdata0(_w_mem_tiles_6_rdata0)
);
M_sprite_layer_mem_tiles_7 __mem__tiles_7(
.clock0(clock),
.clock1(clock),
.in_tiles_7_addr0(_t_tiles_7_addr0),
.in_tiles_7_wenable1(_t_tiles_7_wenable1),
.in_tiles_7_wdata1(_t_tiles_7_wdata1),
.in_tiles_7_addr1(_t_tiles_7_addr1),
.out_tiles_7_rdata0(_w_mem_tiles_7_rdata0)
);
M_sprite_layer_mem_tiles_8 __mem__tiles_8(
.clock0(clock),
.clock1(clock),
.in_tiles_8_addr0(_t_tiles_8_addr0),
.in_tiles_8_wenable1(_t_tiles_8_wenable1),
.in_tiles_8_wdata1(_t_tiles_8_wdata1),
.in_tiles_8_addr1(_t_tiles_8_addr1),
.out_tiles_8_rdata0(_w_mem_tiles_8_rdata0)
);
M_sprite_layer_mem_tiles_9 __mem__tiles_9(
.clock0(clock),
.clock1(clock),
.in_tiles_9_addr0(_t_tiles_9_addr0),
.in_tiles_9_wenable1(_t_tiles_9_wenable1),
.in_tiles_9_wdata1(_t_tiles_9_wdata1),
.in_tiles_9_addr1(_t_tiles_9_addr1),
.out_tiles_9_rdata0(_w_mem_tiles_9_rdata0)
);
M_sprite_layer_mem_tiles_10 __mem__tiles_10(
.clock0(clock),
.clock1(clock),
.in_tiles_10_addr0(_t_tiles_10_addr0),
.in_tiles_10_wenable1(_t_tiles_10_wenable1),
.in_tiles_10_wdata1(_t_tiles_10_wdata1),
.in_tiles_10_addr1(_t_tiles_10_addr1),
.out_tiles_10_rdata0(_w_mem_tiles_10_rdata0)
);
M_sprite_layer_mem_tiles_11 __mem__tiles_11(
.clock0(clock),
.clock1(clock),
.in_tiles_11_addr0(_t_tiles_11_addr0),
.in_tiles_11_wenable1(_t_tiles_11_wenable1),
.in_tiles_11_wdata1(_t_tiles_11_wdata1),
.in_tiles_11_addr1(_t_tiles_11_addr1),
.out_tiles_11_rdata0(_w_mem_tiles_11_rdata0)
);
M_sprite_layer_mem_tiles_12 __mem__tiles_12(
.clock0(clock),
.clock1(clock),
.in_tiles_12_addr0(_t_tiles_12_addr0),
.in_tiles_12_wenable1(_t_tiles_12_wenable1),
.in_tiles_12_wdata1(_t_tiles_12_wdata1),
.in_tiles_12_addr1(_t_tiles_12_addr1),
.out_tiles_12_rdata0(_w_mem_tiles_12_rdata0)
);

assign _w_sprite_to_negative = _q_sprite_double[in_sprite_set_number]?-31:-15;
assign _w_deltax = {{7{in_sprite_update[4+:1]}},in_sprite_update[0+:4]};
assign _w_pix_visible_11 = _d_sprite_active[11]&&_w_xinrange_11&&_w_yinrange_11&&(_w_mem_tiles_11_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[11])>>>_q_sprite_double[11]))+:1]);
assign _w_yinrange_11 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[11]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[11]+_w_spritesize_11));
assign _w_xinrange_11 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[11]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[11]+_w_spritesize_11));
assign _w_pix_visible_10 = _d_sprite_active[10]&&_w_xinrange_10&&_w_yinrange_10&&(_w_mem_tiles_10_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[10])>>>_q_sprite_double[10]))+:1]);
assign _w_yinrange_10 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[10]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[10]+_w_spritesize_10));
assign _w_xinrange_10 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[10]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[10]+_w_spritesize_10));
assign _w_spritesize_9 = _d_sprite_double[9]?32:16;
assign _w_yinrange_12 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[12]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[12]+_w_spritesize_12));
assign _w_yinrange_8 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[8]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[8]+_w_spritesize_8));
assign _w_spritesize_8 = _d_sprite_double[8]?32:16;
assign _w_pix_visible_7 = _d_sprite_active[7]&&_w_xinrange_7&&_w_yinrange_7&&(_w_mem_tiles_7_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[7])>>>_q_sprite_double[7]))+:1]);
assign _w_xinrange_7 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[7]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[7]+_w_spritesize_7));
assign _w_spritesize_3 = _d_sprite_double[3]?32:16;
assign _w_xinrange_9 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[9]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[9]+_w_spritesize_9));
assign _w_yinrange_3 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[3]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[3]+_w_spritesize_3));
assign _w_spritesize_12 = _d_sprite_double[12]?32:16;
assign _w_yinrange_2 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[2]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[2]+_w_spritesize_2));
assign _w_yinrange_6 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[6]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[6]+_w_spritesize_6));
assign _w_pix_visible_2 = _d_sprite_active[2]&&_w_xinrange_2&&_w_yinrange_2&&(_w_mem_tiles_2_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[2])>>>_q_sprite_double[2]))+:1]);
assign _w_sprite_offscreen_x = ($signed(_q_sprite_x[in_sprite_set_number])<$signed(_w_sprite_offscreen_negative))||($signed(_q_sprite_x[in_sprite_set_number])>$signed(640));
assign _w_pix_visible_9 = _d_sprite_active[9]&&_w_xinrange_9&&_w_yinrange_9&&(_w_mem_tiles_9_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[9])>>>_q_sprite_double[9]))+:1]);
assign _w_spritesize_4 = _d_sprite_double[4]?32:16;
assign _w_xinrange_5 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[5]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[5]+_w_spritesize_5));
assign _w_spritesize_5 = _d_sprite_double[5]?32:16;
assign _w_pix_visible_3 = _d_sprite_active[3]&&_w_xinrange_3&&_w_yinrange_3&&(_w_mem_tiles_3_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[3])>>>_q_sprite_double[3]))+:1]);
assign _w_pix_visible_1 = _d_sprite_active[1]&&_w_xinrange_1&&_w_yinrange_1&&(_w_mem_tiles_1_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[1])>>>_q_sprite_double[1]))+:1]);
assign _w_xinrange_2 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[2]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[2]+_w_spritesize_2));
assign _w_sprite_offscreen_negative = _q_sprite_double[in_sprite_set_number]?-32:-16;
assign _w_spritesize_2 = _d_sprite_double[2]?32:16;
assign _w_pix_visible_8 = _d_sprite_active[8]&&_w_xinrange_8&&_w_yinrange_8&&(_w_mem_tiles_8_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[8])>>>_q_sprite_double[8]))+:1]);
assign _w_spritesize_1 = _d_sprite_double[1]?32:16;
assign _w_xinrange_1 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[1]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[1]+_w_spritesize_1));
assign _w_xinrange_8 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[8]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[8]+_w_spritesize_8));
assign _w_pix_visible_0 = _d_sprite_active[0]&&_w_xinrange_0&&_w_yinrange_0&&(_w_mem_tiles_0_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[0])>>>_q_sprite_double[0]))+:1]);
assign _w_spritesize_0 = _d_sprite_double[0]?32:16;
assign _w_pix_visible_12 = _d_sprite_active[12]&&_w_xinrange_12&&_w_yinrange_12&&(_w_mem_tiles_12_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[12])>>>_q_sprite_double[12]))+:1]);
assign _w_xinrange_0 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[0]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[0]+_w_spritesize_0));
assign _w_xinrange_4 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[4]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[4]+_w_spritesize_4));
assign _w_yinrange_1 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[1]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[1]+_w_spritesize_1));
assign _w_yinrange_0 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[0]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[0]+_w_spritesize_0));
assign _w_yinrange_9 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[9]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[9]+_w_spritesize_9));
assign _w_xinrange_3 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[3]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[3]+_w_spritesize_3));
assign _w_sprite_offscreen_y = ($signed(_q_sprite_y[in_sprite_set_number])<$signed(_w_sprite_offscreen_negative))||($signed(_q_sprite_y[in_sprite_set_number])>$signed(480));
assign _w_yinrange_4 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[4]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[4]+_w_spritesize_4));
assign _w_pix_visible_4 = _d_sprite_active[4]&&_w_xinrange_4&&_w_yinrange_4&&(_w_mem_tiles_4_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[4])>>>_q_sprite_double[4]))+:1]);
assign _w_xinrange_12 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[12]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[12]+_w_spritesize_12));
assign _w_spritesize_10 = _d_sprite_double[10]?32:16;
assign _w_yinrange_7 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[7]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[7]+_w_spritesize_7));
assign _w_xinrange_6 = ($signed({1'b0,in_pix_x})>=$signed(_d_sprite_x[6]))&&($signed({1'b0,in_pix_x})<$signed(_d_sprite_x[6]+_w_spritesize_6));
assign _w_yinrange_5 = ($signed({1'b0,in_pix_y})>=$signed(_d_sprite_y[5]))&&($signed({1'b0,in_pix_y})<$signed(_d_sprite_y[5]+_w_spritesize_5));
assign _w_spritesize_11 = _d_sprite_double[11]?32:16;
assign _w_pix_visible_5 = _d_sprite_active[5]&&_w_xinrange_5&&_w_yinrange_5&&(_w_mem_tiles_5_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[5])>>>_q_sprite_double[5]))+:1]);
assign _w_spritesize_6 = _d_sprite_double[6]?32:16;
assign _w_pix_visible_6 = _d_sprite_active[6]&&_w_xinrange_6&&_w_yinrange_6&&(_w_mem_tiles_6_rdata0[(15-(($signed({1'b0,in_pix_x})-_q_sprite_x[6])>>>_q_sprite_double[6]))+:1]);
assign _w_deltay = {{7{in_sprite_update[9+:1]}},in_sprite_update[5+:4]};
assign _w_spritesize_7 = _d_sprite_double[7]?32:16;

always @* begin
_d_sprite_active[0] = _q_sprite_active[0];
_d_sprite_active[1] = _q_sprite_active[1];
_d_sprite_active[2] = _q_sprite_active[2];
_d_sprite_active[3] = _q_sprite_active[3];
_d_sprite_active[4] = _q_sprite_active[4];
_d_sprite_active[5] = _q_sprite_active[5];
_d_sprite_active[6] = _q_sprite_active[6];
_d_sprite_active[7] = _q_sprite_active[7];
_d_sprite_active[8] = _q_sprite_active[8];
_d_sprite_active[9] = _q_sprite_active[9];
_d_sprite_active[10] = _q_sprite_active[10];
_d_sprite_active[11] = _q_sprite_active[11];
_d_sprite_active[12] = _q_sprite_active[12];
_d_sprite_double[0] = _q_sprite_double[0];
_d_sprite_double[1] = _q_sprite_double[1];
_d_sprite_double[2] = _q_sprite_double[2];
_d_sprite_double[3] = _q_sprite_double[3];
_d_sprite_double[4] = _q_sprite_double[4];
_d_sprite_double[5] = _q_sprite_double[5];
_d_sprite_double[6] = _q_sprite_double[6];
_d_sprite_double[7] = _q_sprite_double[7];
_d_sprite_double[8] = _q_sprite_double[8];
_d_sprite_double[9] = _q_sprite_double[9];
_d_sprite_double[10] = _q_sprite_double[10];
_d_sprite_double[11] = _q_sprite_double[11];
_d_sprite_double[12] = _q_sprite_double[12];
_d_sprite_x[0] = _q_sprite_x[0];
_d_sprite_x[1] = _q_sprite_x[1];
_d_sprite_x[2] = _q_sprite_x[2];
_d_sprite_x[3] = _q_sprite_x[3];
_d_sprite_x[4] = _q_sprite_x[4];
_d_sprite_x[5] = _q_sprite_x[5];
_d_sprite_x[6] = _q_sprite_x[6];
_d_sprite_x[7] = _q_sprite_x[7];
_d_sprite_x[8] = _q_sprite_x[8];
_d_sprite_x[9] = _q_sprite_x[9];
_d_sprite_x[10] = _q_sprite_x[10];
_d_sprite_x[11] = _q_sprite_x[11];
_d_sprite_x[12] = _q_sprite_x[12];
_d_sprite_y[0] = _q_sprite_y[0];
_d_sprite_y[1] = _q_sprite_y[1];
_d_sprite_y[2] = _q_sprite_y[2];
_d_sprite_y[3] = _q_sprite_y[3];
_d_sprite_y[4] = _q_sprite_y[4];
_d_sprite_y[5] = _q_sprite_y[5];
_d_sprite_y[6] = _q_sprite_y[6];
_d_sprite_y[7] = _q_sprite_y[7];
_d_sprite_y[8] = _q_sprite_y[8];
_d_sprite_y[9] = _q_sprite_y[9];
_d_sprite_y[10] = _q_sprite_y[10];
_d_sprite_y[11] = _q_sprite_y[11];
_d_sprite_y[12] = _q_sprite_y[12];
_d_sprite_colour[0] = _q_sprite_colour[0];
_d_sprite_colour[1] = _q_sprite_colour[1];
_d_sprite_colour[2] = _q_sprite_colour[2];
_d_sprite_colour[3] = _q_sprite_colour[3];
_d_sprite_colour[4] = _q_sprite_colour[4];
_d_sprite_colour[5] = _q_sprite_colour[5];
_d_sprite_colour[6] = _q_sprite_colour[6];
_d_sprite_colour[7] = _q_sprite_colour[7];
_d_sprite_colour[8] = _q_sprite_colour[8];
_d_sprite_colour[9] = _q_sprite_colour[9];
_d_sprite_colour[10] = _q_sprite_colour[10];
_d_sprite_colour[11] = _q_sprite_colour[11];
_d_sprite_colour[12] = _q_sprite_colour[12];
_d_sprite_tile_number[0] = _q_sprite_tile_number[0];
_d_sprite_tile_number[1] = _q_sprite_tile_number[1];
_d_sprite_tile_number[2] = _q_sprite_tile_number[2];
_d_sprite_tile_number[3] = _q_sprite_tile_number[3];
_d_sprite_tile_number[4] = _q_sprite_tile_number[4];
_d_sprite_tile_number[5] = _q_sprite_tile_number[5];
_d_sprite_tile_number[6] = _q_sprite_tile_number[6];
_d_sprite_tile_number[7] = _q_sprite_tile_number[7];
_d_sprite_tile_number[8] = _q_sprite_tile_number[8];
_d_sprite_tile_number[9] = _q_sprite_tile_number[9];
_d_sprite_tile_number[10] = _q_sprite_tile_number[10];
_d_sprite_tile_number[11] = _q_sprite_tile_number[11];
_d_sprite_tile_number[12] = _q_sprite_tile_number[12];
_d_output_collisions = _q_output_collisions;
_d_detect_collision_0 = _q_detect_collision_0;
_d_detect_collision_1 = _q_detect_collision_1;
_d_detect_collision_2 = _q_detect_collision_2;
_d_detect_collision_3 = _q_detect_collision_3;
_d_detect_collision_4 = _q_detect_collision_4;
_d_detect_collision_5 = _q_detect_collision_5;
_d_detect_collision_6 = _q_detect_collision_6;
_d_detect_collision_7 = _q_detect_collision_7;
_d_detect_collision_8 = _q_detect_collision_8;
_d_detect_collision_9 = _q_detect_collision_9;
_d_detect_collision_10 = _q_detect_collision_10;
_d_detect_collision_11 = _q_detect_collision_11;
_d_detect_collision_12 = _q_detect_collision_12;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_sprite_layer_display = _q_sprite_layer_display;
_d_sprite_read_active = _q_sprite_read_active;
_d_sprite_read_double = _q_sprite_read_double;
_d_sprite_read_colour = _q_sprite_read_colour;
_d_sprite_read_x = _q_sprite_read_x;
_d_sprite_read_y = _q_sprite_read_y;
_d_sprite_read_tile = _q_sprite_read_tile;
_d_collision_0 = _q_collision_0;
_d_collision_1 = _q_collision_1;
_d_collision_2 = _q_collision_2;
_d_collision_3 = _q_collision_3;
_d_collision_4 = _q_collision_4;
_d_collision_5 = _q_collision_5;
_d_collision_6 = _q_collision_6;
_d_collision_7 = _q_collision_7;
_d_collision_8 = _q_collision_8;
_d_collision_9 = _q_collision_9;
_d_collision_10 = _q_collision_10;
_d_collision_11 = _q_collision_11;
_d_collision_12 = _q_collision_12;
_d_index = _q_index;
_t_tiles_0_addr0 = 0;
_t_tiles_0_wenable1 = 0;
_t_tiles_0_wdata1 = 0;
_t_tiles_0_addr1 = 0;
_t_tiles_1_addr0 = 0;
_t_tiles_1_wenable1 = 0;
_t_tiles_1_wdata1 = 0;
_t_tiles_1_addr1 = 0;
_t_tiles_2_addr0 = 0;
_t_tiles_2_wenable1 = 0;
_t_tiles_2_wdata1 = 0;
_t_tiles_2_addr1 = 0;
_t_tiles_3_addr0 = 0;
_t_tiles_3_wenable1 = 0;
_t_tiles_3_wdata1 = 0;
_t_tiles_3_addr1 = 0;
_t_tiles_4_addr0 = 0;
_t_tiles_4_wenable1 = 0;
_t_tiles_4_wdata1 = 0;
_t_tiles_4_addr1 = 0;
_t_tiles_5_addr0 = 0;
_t_tiles_5_wenable1 = 0;
_t_tiles_5_wdata1 = 0;
_t_tiles_5_addr1 = 0;
_t_tiles_6_addr0 = 0;
_t_tiles_6_wenable1 = 0;
_t_tiles_6_wdata1 = 0;
_t_tiles_6_addr1 = 0;
_t_tiles_7_addr0 = 0;
_t_tiles_7_wenable1 = 0;
_t_tiles_7_wdata1 = 0;
_t_tiles_7_addr1 = 0;
_t_tiles_8_addr0 = 0;
_t_tiles_8_wenable1 = 0;
_t_tiles_8_wdata1 = 0;
_t_tiles_8_addr1 = 0;
_t_tiles_9_addr0 = 0;
_t_tiles_9_wenable1 = 0;
_t_tiles_9_wdata1 = 0;
_t_tiles_9_addr1 = 0;
_t_tiles_10_addr0 = 0;
_t_tiles_10_wenable1 = 0;
_t_tiles_10_wdata1 = 0;
_t_tiles_10_addr1 = 0;
_t_tiles_11_addr0 = 0;
_t_tiles_11_wenable1 = 0;
_t_tiles_11_wdata1 = 0;
_t_tiles_11_addr1 = 0;
_t_tiles_12_addr0 = 0;
_t_tiles_12_wenable1 = 0;
_t_tiles_12_wdata1 = 0;
_t_tiles_12_addr1 = 0;
// _always_pre
_t_tiles_0_addr0 = _q_sprite_tile_number[0]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[0])>>>_q_sprite_double[0]);
_t_tiles_0_wenable1 = 1;
_d_collision_0 = (_q_output_collisions)?_q_detect_collision_0:_q_collision_0;
_t_tiles_1_addr0 = _q_sprite_tile_number[1]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[1])>>>_q_sprite_double[1]);
_t_tiles_1_wenable1 = 1;
_d_collision_1 = (_q_output_collisions)?_q_detect_collision_1:_q_collision_1;
_t_tiles_2_addr0 = _q_sprite_tile_number[2]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[2])>>>_q_sprite_double[2]);
_t_tiles_2_wenable1 = 1;
_d_collision_2 = (_q_output_collisions)?_q_detect_collision_2:_q_collision_2;
_t_tiles_3_addr0 = _q_sprite_tile_number[3]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[3])>>>_q_sprite_double[3]);
_t_tiles_3_wenable1 = 1;
_d_collision_3 = (_q_output_collisions)?_q_detect_collision_3:_q_collision_3;
_t_tiles_4_addr0 = _q_sprite_tile_number[4]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[4])>>>_q_sprite_double[4]);
_t_tiles_4_wenable1 = 1;
_d_collision_4 = (_q_output_collisions)?_q_detect_collision_4:_q_collision_4;
_t_tiles_5_addr0 = _q_sprite_tile_number[5]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[5])>>>_q_sprite_double[5]);
_t_tiles_5_wenable1 = 1;
_d_collision_5 = (_q_output_collisions)?_q_detect_collision_5:_q_collision_5;
_t_tiles_6_addr0 = _q_sprite_tile_number[6]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[6])>>>_q_sprite_double[6]);
_t_tiles_6_wenable1 = 1;
_d_collision_6 = (_q_output_collisions)?_q_detect_collision_6:_q_collision_6;
_t_tiles_7_addr0 = _q_sprite_tile_number[7]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[7])>>>_q_sprite_double[7]);
_t_tiles_7_wenable1 = 1;
_d_collision_7 = (_q_output_collisions)?_q_detect_collision_7:_q_collision_7;
_t_tiles_8_addr0 = _q_sprite_tile_number[8]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[8])>>>_q_sprite_double[8]);
_t_tiles_8_wenable1 = 1;
_d_collision_8 = (_q_output_collisions)?_q_detect_collision_8:_q_collision_8;
_t_tiles_9_addr0 = _q_sprite_tile_number[9]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[9])>>>_q_sprite_double[9]);
_t_tiles_9_wenable1 = 1;
_d_collision_9 = (_q_output_collisions)?_q_detect_collision_9:_q_collision_9;
_t_tiles_10_addr0 = _q_sprite_tile_number[10]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[10])>>>_q_sprite_double[10]);
_t_tiles_10_wenable1 = 1;
_d_collision_10 = (_q_output_collisions)?_q_detect_collision_10:_q_collision_10;
_t_tiles_11_addr0 = _q_sprite_tile_number[11]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[11])>>>_q_sprite_double[11]);
_t_tiles_11_wenable1 = 1;
_d_collision_11 = (_q_output_collisions)?_q_detect_collision_11:_q_collision_11;
_t_tiles_12_addr0 = _q_sprite_tile_number[12]*16+(($signed({1'b0,in_pix_y})-_q_sprite_y[12])>>>_q_sprite_double[12]);
_t_tiles_12_wenable1 = 1;
_d_collision_12 = (_q_output_collisions)?_q_detect_collision_12:_q_collision_12;
_d_sprite_layer_display = 0;
_d_sprite_read_active = _q_sprite_active[in_sprite_set_number];
_d_sprite_read_double = _q_sprite_double[in_sprite_set_number];
_d_sprite_read_colour = _q_sprite_colour[in_sprite_set_number];
_d_sprite_read_x = _q_sprite_x[in_sprite_set_number];
_d_sprite_read_y = _q_sprite_y[in_sprite_set_number];
_d_sprite_read_tile = _q_sprite_tile_number[in_sprite_set_number];
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_output_collisions = 0;
_t_tiles_0_addr0 = 0;
_t_tiles_0_wenable1 = 0;
_t_tiles_0_wdata1 = 0;
_t_tiles_0_addr1 = 0;
_t_tiles_1_addr0 = 0;
_t_tiles_1_wenable1 = 0;
_t_tiles_1_wdata1 = 0;
_t_tiles_1_addr1 = 0;
_t_tiles_2_addr0 = 0;
_t_tiles_2_wenable1 = 0;
_t_tiles_2_wdata1 = 0;
_t_tiles_2_addr1 = 0;
_t_tiles_3_addr0 = 0;
_t_tiles_3_wenable1 = 0;
_t_tiles_3_wdata1 = 0;
_t_tiles_3_addr1 = 0;
_t_tiles_4_addr0 = 0;
_t_tiles_4_wenable1 = 0;
_t_tiles_4_wdata1 = 0;
_t_tiles_4_addr1 = 0;
_t_tiles_5_addr0 = 0;
_t_tiles_5_wenable1 = 0;
_t_tiles_5_wdata1 = 0;
_t_tiles_5_addr1 = 0;
_t_tiles_6_addr0 = 0;
_t_tiles_6_wenable1 = 0;
_t_tiles_6_wdata1 = 0;
_t_tiles_6_addr1 = 0;
_t_tiles_7_addr0 = 0;
_t_tiles_7_wenable1 = 0;
_t_tiles_7_wdata1 = 0;
_t_tiles_7_addr1 = 0;
_t_tiles_8_addr0 = 0;
_t_tiles_8_wenable1 = 0;
_t_tiles_8_wdata1 = 0;
_t_tiles_8_addr1 = 0;
_t_tiles_9_addr0 = 0;
_t_tiles_9_wenable1 = 0;
_t_tiles_9_wdata1 = 0;
_t_tiles_9_addr1 = 0;
_t_tiles_10_addr0 = 0;
_t_tiles_10_wenable1 = 0;
_t_tiles_10_wdata1 = 0;
_t_tiles_10_addr1 = 0;
_t_tiles_11_addr0 = 0;
_t_tiles_11_wenable1 = 0;
_t_tiles_11_wdata1 = 0;
_t_tiles_11_addr1 = 0;
_t_tiles_12_addr0 = 0;
_t_tiles_12_wenable1 = 0;
_t_tiles_12_wdata1 = 0;
_t_tiles_12_addr1 = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_pix_vblank) begin
// __block_5
// __block_7
if (~_q_output_collisions) begin
// __block_8
// __block_10
_d_detect_collision_0 = 0;
_d_detect_collision_1 = 0;
_d_detect_collision_2 = 0;
_d_detect_collision_3 = 0;
_d_detect_collision_4 = 0;
_d_detect_collision_5 = 0;
_d_detect_collision_6 = 0;
_d_detect_collision_7 = 0;
_d_detect_collision_8 = 0;
_d_detect_collision_9 = 0;
_d_detect_collision_10 = 0;
_d_detect_collision_11 = 0;
_d_detect_collision_12 = 0;
// __block_11
end else begin
// __block_9
// __block_12
_d_output_collisions = 0;
// __block_13
end
// __block_14
// __block_15
end else begin
// __block_6
// __block_16
if (in_pix_active) begin
// __block_17
// __block_19
if ((_w_pix_visible_0)) begin
// __block_20
// __block_22
_d_pix_red = _q_sprite_colour[0][4+:2];
_d_pix_green = _q_sprite_colour[0][2+:2];
_d_pix_blue = _q_sprite_colour[0][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_0 = _q_detect_collision_0|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_23
end else begin
// __block_21
end
// __block_24
if ((_w_pix_visible_1)) begin
// __block_25
// __block_27
_d_pix_red = _q_sprite_colour[1][4+:2];
_d_pix_green = _q_sprite_colour[1][2+:2];
_d_pix_blue = _q_sprite_colour[1][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_1 = _q_detect_collision_1|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_28
end else begin
// __block_26
end
// __block_29
if ((_w_pix_visible_2)) begin
// __block_30
// __block_32
_d_pix_red = _q_sprite_colour[2][4+:2];
_d_pix_green = _q_sprite_colour[2][2+:2];
_d_pix_blue = _q_sprite_colour[2][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_2 = _q_detect_collision_2|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_33
end else begin
// __block_31
end
// __block_34
if ((_w_pix_visible_3)) begin
// __block_35
// __block_37
_d_pix_red = _q_sprite_colour[3][4+:2];
_d_pix_green = _q_sprite_colour[3][2+:2];
_d_pix_blue = _q_sprite_colour[3][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_3 = _q_detect_collision_3|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_38
end else begin
// __block_36
end
// __block_39
if ((_w_pix_visible_4)) begin
// __block_40
// __block_42
_d_pix_red = _q_sprite_colour[4][4+:2];
_d_pix_green = _q_sprite_colour[4][2+:2];
_d_pix_blue = _q_sprite_colour[4][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_4 = _q_detect_collision_4|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_43
end else begin
// __block_41
end
// __block_44
if ((_w_pix_visible_5)) begin
// __block_45
// __block_47
_d_pix_red = _q_sprite_colour[5][4+:2];
_d_pix_green = _q_sprite_colour[5][2+:2];
_d_pix_blue = _q_sprite_colour[5][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_5 = _q_detect_collision_5|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_48
end else begin
// __block_46
end
// __block_49
if ((_w_pix_visible_6)) begin
// __block_50
// __block_52
_d_pix_red = _q_sprite_colour[6][4+:2];
_d_pix_green = _q_sprite_colour[6][2+:2];
_d_pix_blue = _q_sprite_colour[6][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_6 = _q_detect_collision_6|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_53
end else begin
// __block_51
end
// __block_54
if ((_w_pix_visible_7)) begin
// __block_55
// __block_57
_d_pix_red = _q_sprite_colour[7][4+:2];
_d_pix_green = _q_sprite_colour[7][2+:2];
_d_pix_blue = _q_sprite_colour[7][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_7 = _q_detect_collision_7|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_58
end else begin
// __block_56
end
// __block_59
if ((_w_pix_visible_8)) begin
// __block_60
// __block_62
_d_pix_red = _q_sprite_colour[8][4+:2];
_d_pix_green = _q_sprite_colour[8][2+:2];
_d_pix_blue = _q_sprite_colour[8][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_8 = _q_detect_collision_8|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_63
end else begin
// __block_61
end
// __block_64
if ((_w_pix_visible_9)) begin
// __block_65
// __block_67
_d_pix_red = _q_sprite_colour[9][4+:2];
_d_pix_green = _q_sprite_colour[9][2+:2];
_d_pix_blue = _q_sprite_colour[9][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_9 = _q_detect_collision_9|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_68
end else begin
// __block_66
end
// __block_69
if ((_w_pix_visible_10)) begin
// __block_70
// __block_72
_d_pix_red = _q_sprite_colour[10][4+:2];
_d_pix_green = _q_sprite_colour[10][2+:2];
_d_pix_blue = _q_sprite_colour[10][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_10 = _q_detect_collision_10|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_73
end else begin
// __block_71
end
// __block_74
if ((_w_pix_visible_11)) begin
// __block_75
// __block_77
_d_pix_red = _q_sprite_colour[11][4+:2];
_d_pix_green = _q_sprite_colour[11][2+:2];
_d_pix_blue = _q_sprite_colour[11][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_11 = _q_detect_collision_11|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_78
end else begin
// __block_76
end
// __block_79
if ((_w_pix_visible_12)) begin
// __block_80
// __block_82
_d_pix_red = _q_sprite_colour[12][4+:2];
_d_pix_green = _q_sprite_colour[12][2+:2];
_d_pix_blue = _q_sprite_colour[12][0+:2];
_d_sprite_layer_display = 1;
_d_detect_collision_12 = _q_detect_collision_12|{in_collision_layer_1,in_collision_layer_2,in_collision_layer_3,_w_pix_visible_12,_w_pix_visible_11,_w_pix_visible_10,_w_pix_visible_9,_w_pix_visible_8,_w_pix_visible_7,_w_pix_visible_6,_w_pix_visible_5,_w_pix_visible_4,_w_pix_visible_3,_w_pix_visible_2,_w_pix_visible_1,_w_pix_visible_0};
// __block_83
end else begin
// __block_81
end
// __block_84
_d_output_collisions = (in_pix_x==639)&&(in_pix_y==479);
// __block_85
end else begin
// __block_18
end
// __block_86
// __block_87
end
// __block_88
if (in_sprite_writer_active) begin
// __block_89
// __block_91
  case (in_sprite_writer_sprite)
  0: begin
// __block_93_case
// __block_94
_t_tiles_0_addr1 = in_sprite_writer_line;
_t_tiles_0_wdata1 = in_sprite_writer_bitmap;
// __block_95
  end
  1: begin
// __block_96_case
// __block_97
_t_tiles_1_addr1 = in_sprite_writer_line;
_t_tiles_1_wdata1 = in_sprite_writer_bitmap;
// __block_98
  end
  2: begin
// __block_99_case
// __block_100
_t_tiles_2_addr1 = in_sprite_writer_line;
_t_tiles_2_wdata1 = in_sprite_writer_bitmap;
// __block_101
  end
  3: begin
// __block_102_case
// __block_103
_t_tiles_3_addr1 = in_sprite_writer_line;
_t_tiles_3_wdata1 = in_sprite_writer_bitmap;
// __block_104
  end
  4: begin
// __block_105_case
// __block_106
_t_tiles_4_addr1 = in_sprite_writer_line;
_t_tiles_4_wdata1 = in_sprite_writer_bitmap;
// __block_107
  end
  5: begin
// __block_108_case
// __block_109
_t_tiles_5_addr1 = in_sprite_writer_line;
_t_tiles_5_wdata1 = in_sprite_writer_bitmap;
// __block_110
  end
  6: begin
// __block_111_case
// __block_112
_t_tiles_6_addr1 = in_sprite_writer_line;
_t_tiles_6_wdata1 = in_sprite_writer_bitmap;
// __block_113
  end
  7: begin
// __block_114_case
// __block_115
_t_tiles_7_addr1 = in_sprite_writer_line;
_t_tiles_7_wdata1 = in_sprite_writer_bitmap;
// __block_116
  end
  8: begin
// __block_117_case
// __block_118
_t_tiles_8_addr1 = in_sprite_writer_line;
_t_tiles_8_wdata1 = in_sprite_writer_bitmap;
// __block_119
  end
  9: begin
// __block_120_case
// __block_121
_t_tiles_9_addr1 = in_sprite_writer_line;
_t_tiles_9_wdata1 = in_sprite_writer_bitmap;
// __block_122
  end
  10: begin
// __block_123_case
// __block_124
_t_tiles_10_addr1 = in_sprite_writer_line;
_t_tiles_10_wdata1 = in_sprite_writer_bitmap;
// __block_125
  end
  11: begin
// __block_126_case
// __block_127
_t_tiles_11_addr1 = in_sprite_writer_line;
_t_tiles_11_wdata1 = in_sprite_writer_bitmap;
// __block_128
  end
  12: begin
// __block_129_case
// __block_130
_t_tiles_12_addr1 = in_sprite_writer_line;
_t_tiles_12_wdata1 = in_sprite_writer_bitmap;
// __block_131
  end
endcase
// __block_92
// __block_132
end else begin
// __block_90
end
// __block_133
  case (in_sprite_layer_write)
  1: begin
// __block_135_case
// __block_136
_d_sprite_active[in_sprite_set_number] = in_sprite_set_active;
// __block_137
  end
  2: begin
// __block_138_case
// __block_139
_d_sprite_tile_number[in_sprite_set_number] = in_sprite_set_tile;
// __block_140
  end
  3: begin
// __block_141_case
// __block_142
_d_sprite_colour[in_sprite_set_number] = in_sprite_set_colour;
// __block_143
  end
  4: begin
// __block_144_case
// __block_145
_d_sprite_x[in_sprite_set_number] = in_sprite_set_x;
// __block_146
  end
  5: begin
// __block_147_case
// __block_148
_d_sprite_y[in_sprite_set_number] = in_sprite_set_y;
// __block_149
  end
  6: begin
// __block_150_case
// __block_151
_d_sprite_double[in_sprite_set_number] = in_sprite_set_double;
// __block_152
  end
  10: begin
// __block_153_case
// __block_154
if (in_sprite_update[10+:1]) begin
// __block_155
// __block_157
_d_sprite_tile_number[in_sprite_set_number] = _q_sprite_tile_number[in_sprite_set_number]+1;
// __block_158
end else begin
// __block_156
end
// __block_159
if (in_sprite_update[11+:1]||in_sprite_update[12+:1]) begin
// __block_160
// __block_162
_d_sprite_active[in_sprite_set_number] = (_w_sprite_offscreen_x||_w_sprite_offscreen_y)?0:_q_sprite_active[in_sprite_set_number];
// __block_163
end else begin
// __block_161
end
// __block_164
_d_sprite_x[in_sprite_set_number] = _w_sprite_offscreen_x?(($signed(_q_sprite_x[in_sprite_set_number])<$signed(_w_sprite_offscreen_negative))?$signed(640):_w_sprite_to_negative):_q_sprite_x[in_sprite_set_number]+_w_deltax;
_d_sprite_y[in_sprite_set_number] = _w_sprite_offscreen_y?(($signed(_q_sprite_y[in_sprite_set_number])<$signed(_w_sprite_offscreen_negative))?$signed(480):_w_sprite_to_negative):_q_sprite_y[in_sprite_set_number]+_w_deltay;
// __block_165
  end
endcase
// __block_134
// __block_166
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of sprite_layer
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_tilemap_mem_tiles16x16(
input      [8:0]                in_tiles16x16_addr0,
output reg  [15:0]     out_tiles16x16_rdata0,
output reg  [15:0]     out_tiles16x16_rdata1,
input      [0:0]             in_tiles16x16_wenable1,
input      [15:0]                 in_tiles16x16_wdata1,
input      [8:0]                in_tiles16x16_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[511:0];
always @(posedge clock0) begin
  out_tiles16x16_rdata0 <= buffer[in_tiles16x16_addr0];
end
always @(posedge clock1) begin
  if (in_tiles16x16_wenable1) begin
    buffer[in_tiles16x16_addr1] <= in_tiles16x16_wdata1;
  end
end
initial begin
 buffer[0] = 0;
 buffer[1] = 0;
 buffer[2] = 0;
 buffer[3] = 0;
 buffer[4] = 0;
 buffer[5] = 0;
 buffer[6] = 0;
 buffer[7] = 0;
 buffer[8] = 0;
 buffer[9] = 0;
 buffer[10] = 0;
 buffer[11] = 0;
 buffer[12] = 0;
 buffer[13] = 0;
 buffer[14] = 0;
 buffer[15] = 0;
 buffer[16] = 0;
 buffer[17] = 0;
 buffer[18] = 0;
 buffer[19] = 0;
 buffer[20] = 0;
 buffer[21] = 0;
 buffer[22] = 0;
 buffer[23] = 0;
 buffer[24] = 0;
 buffer[25] = 0;
 buffer[26] = 0;
 buffer[27] = 0;
 buffer[28] = 0;
 buffer[29] = 0;
 buffer[30] = 0;
 buffer[31] = 0;
 buffer[32] = 0;
 buffer[33] = 0;
 buffer[34] = 0;
 buffer[35] = 0;
 buffer[36] = 0;
 buffer[37] = 0;
 buffer[38] = 0;
 buffer[39] = 0;
 buffer[40] = 0;
 buffer[41] = 0;
 buffer[42] = 0;
 buffer[43] = 0;
 buffer[44] = 0;
 buffer[45] = 0;
 buffer[46] = 0;
 buffer[47] = 0;
 buffer[48] = 0;
 buffer[49] = 0;
 buffer[50] = 0;
 buffer[51] = 0;
 buffer[52] = 0;
 buffer[53] = 0;
 buffer[54] = 0;
 buffer[55] = 0;
 buffer[56] = 0;
 buffer[57] = 0;
 buffer[58] = 0;
 buffer[59] = 0;
 buffer[60] = 0;
 buffer[61] = 0;
 buffer[62] = 0;
 buffer[63] = 0;
 buffer[64] = 0;
 buffer[65] = 0;
 buffer[66] = 0;
 buffer[67] = 0;
 buffer[68] = 0;
 buffer[69] = 0;
 buffer[70] = 0;
 buffer[71] = 0;
 buffer[72] = 0;
 buffer[73] = 0;
 buffer[74] = 0;
 buffer[75] = 0;
 buffer[76] = 0;
 buffer[77] = 0;
 buffer[78] = 0;
 buffer[79] = 0;
 buffer[80] = 0;
 buffer[81] = 0;
 buffer[82] = 0;
 buffer[83] = 0;
 buffer[84] = 0;
 buffer[85] = 0;
 buffer[86] = 0;
 buffer[87] = 0;
 buffer[88] = 0;
 buffer[89] = 0;
 buffer[90] = 0;
 buffer[91] = 0;
 buffer[92] = 0;
 buffer[93] = 0;
 buffer[94] = 0;
 buffer[95] = 0;
 buffer[96] = 0;
 buffer[97] = 0;
 buffer[98] = 0;
 buffer[99] = 0;
 buffer[100] = 0;
 buffer[101] = 0;
 buffer[102] = 0;
 buffer[103] = 0;
 buffer[104] = 0;
 buffer[105] = 0;
 buffer[106] = 0;
 buffer[107] = 0;
 buffer[108] = 0;
 buffer[109] = 0;
 buffer[110] = 0;
 buffer[111] = 0;
 buffer[112] = 0;
 buffer[113] = 0;
 buffer[114] = 0;
 buffer[115] = 0;
 buffer[116] = 0;
 buffer[117] = 0;
 buffer[118] = 0;
 buffer[119] = 0;
 buffer[120] = 0;
 buffer[121] = 0;
 buffer[122] = 0;
 buffer[123] = 0;
 buffer[124] = 0;
 buffer[125] = 0;
 buffer[126] = 0;
 buffer[127] = 0;
 buffer[128] = 0;
 buffer[129] = 0;
 buffer[130] = 0;
 buffer[131] = 0;
 buffer[132] = 0;
 buffer[133] = 0;
 buffer[134] = 0;
 buffer[135] = 0;
 buffer[136] = 0;
 buffer[137] = 0;
 buffer[138] = 0;
 buffer[139] = 0;
 buffer[140] = 0;
 buffer[141] = 0;
 buffer[142] = 0;
 buffer[143] = 0;
 buffer[144] = 0;
 buffer[145] = 0;
 buffer[146] = 0;
 buffer[147] = 0;
 buffer[148] = 0;
 buffer[149] = 0;
 buffer[150] = 0;
 buffer[151] = 0;
 buffer[152] = 0;
 buffer[153] = 0;
 buffer[154] = 0;
 buffer[155] = 0;
 buffer[156] = 0;
 buffer[157] = 0;
 buffer[158] = 0;
 buffer[159] = 0;
 buffer[160] = 0;
 buffer[161] = 0;
 buffer[162] = 0;
 buffer[163] = 0;
 buffer[164] = 0;
 buffer[165] = 0;
 buffer[166] = 0;
 buffer[167] = 0;
 buffer[168] = 0;
 buffer[169] = 0;
 buffer[170] = 0;
 buffer[171] = 0;
 buffer[172] = 0;
 buffer[173] = 0;
 buffer[174] = 0;
 buffer[175] = 0;
 buffer[176] = 0;
 buffer[177] = 0;
 buffer[178] = 0;
 buffer[179] = 0;
 buffer[180] = 0;
 buffer[181] = 0;
 buffer[182] = 0;
 buffer[183] = 0;
 buffer[184] = 0;
 buffer[185] = 0;
 buffer[186] = 0;
 buffer[187] = 0;
 buffer[188] = 0;
 buffer[189] = 0;
 buffer[190] = 0;
 buffer[191] = 0;
 buffer[192] = 0;
 buffer[193] = 0;
 buffer[194] = 0;
 buffer[195] = 0;
 buffer[196] = 0;
 buffer[197] = 0;
 buffer[198] = 0;
 buffer[199] = 0;
 buffer[200] = 0;
 buffer[201] = 0;
 buffer[202] = 0;
 buffer[203] = 0;
 buffer[204] = 0;
 buffer[205] = 0;
 buffer[206] = 0;
 buffer[207] = 0;
 buffer[208] = 0;
 buffer[209] = 0;
 buffer[210] = 0;
 buffer[211] = 0;
 buffer[212] = 0;
 buffer[213] = 0;
 buffer[214] = 0;
 buffer[215] = 0;
 buffer[216] = 0;
 buffer[217] = 0;
 buffer[218] = 0;
 buffer[219] = 0;
 buffer[220] = 0;
 buffer[221] = 0;
 buffer[222] = 0;
 buffer[223] = 0;
 buffer[224] = 0;
 buffer[225] = 0;
 buffer[226] = 0;
 buffer[227] = 0;
 buffer[228] = 0;
 buffer[229] = 0;
 buffer[230] = 0;
 buffer[231] = 0;
 buffer[232] = 0;
 buffer[233] = 0;
 buffer[234] = 0;
 buffer[235] = 0;
 buffer[236] = 0;
 buffer[237] = 0;
 buffer[238] = 0;
 buffer[239] = 0;
 buffer[240] = 0;
 buffer[241] = 0;
 buffer[242] = 0;
 buffer[243] = 0;
 buffer[244] = 0;
 buffer[245] = 0;
 buffer[246] = 0;
 buffer[247] = 0;
 buffer[248] = 0;
 buffer[249] = 0;
 buffer[250] = 0;
 buffer[251] = 0;
 buffer[252] = 0;
 buffer[253] = 0;
 buffer[254] = 0;
 buffer[255] = 0;
 buffer[256] = 0;
 buffer[257] = 0;
 buffer[258] = 0;
 buffer[259] = 0;
 buffer[260] = 0;
 buffer[261] = 0;
 buffer[262] = 0;
 buffer[263] = 0;
 buffer[264] = 0;
 buffer[265] = 0;
 buffer[266] = 0;
 buffer[267] = 0;
 buffer[268] = 0;
 buffer[269] = 0;
 buffer[270] = 0;
 buffer[271] = 0;
 buffer[272] = 0;
 buffer[273] = 0;
 buffer[274] = 0;
 buffer[275] = 0;
 buffer[276] = 0;
 buffer[277] = 0;
 buffer[278] = 0;
 buffer[279] = 0;
 buffer[280] = 0;
 buffer[281] = 0;
 buffer[282] = 0;
 buffer[283] = 0;
 buffer[284] = 0;
 buffer[285] = 0;
 buffer[286] = 0;
 buffer[287] = 0;
 buffer[288] = 0;
 buffer[289] = 0;
 buffer[290] = 0;
 buffer[291] = 0;
 buffer[292] = 0;
 buffer[293] = 0;
 buffer[294] = 0;
 buffer[295] = 0;
 buffer[296] = 0;
 buffer[297] = 0;
 buffer[298] = 0;
 buffer[299] = 0;
 buffer[300] = 0;
 buffer[301] = 0;
 buffer[302] = 0;
 buffer[303] = 0;
 buffer[304] = 0;
 buffer[305] = 0;
 buffer[306] = 0;
 buffer[307] = 0;
 buffer[308] = 0;
 buffer[309] = 0;
 buffer[310] = 0;
 buffer[311] = 0;
 buffer[312] = 0;
 buffer[313] = 0;
 buffer[314] = 0;
 buffer[315] = 0;
 buffer[316] = 0;
 buffer[317] = 0;
 buffer[318] = 0;
 buffer[319] = 0;
 buffer[320] = 0;
 buffer[321] = 0;
 buffer[322] = 0;
 buffer[323] = 0;
 buffer[324] = 0;
 buffer[325] = 0;
 buffer[326] = 0;
 buffer[327] = 0;
 buffer[328] = 0;
 buffer[329] = 0;
 buffer[330] = 0;
 buffer[331] = 0;
 buffer[332] = 0;
 buffer[333] = 0;
 buffer[334] = 0;
 buffer[335] = 0;
 buffer[336] = 0;
 buffer[337] = 0;
 buffer[338] = 0;
 buffer[339] = 0;
 buffer[340] = 0;
 buffer[341] = 0;
 buffer[342] = 0;
 buffer[343] = 0;
 buffer[344] = 0;
 buffer[345] = 0;
 buffer[346] = 0;
 buffer[347] = 0;
 buffer[348] = 0;
 buffer[349] = 0;
 buffer[350] = 0;
 buffer[351] = 0;
 buffer[352] = 0;
 buffer[353] = 0;
 buffer[354] = 0;
 buffer[355] = 0;
 buffer[356] = 0;
 buffer[357] = 0;
 buffer[358] = 0;
 buffer[359] = 0;
 buffer[360] = 0;
 buffer[361] = 0;
 buffer[362] = 0;
 buffer[363] = 0;
 buffer[364] = 0;
 buffer[365] = 0;
 buffer[366] = 0;
 buffer[367] = 0;
 buffer[368] = 0;
 buffer[369] = 0;
 buffer[370] = 0;
 buffer[371] = 0;
 buffer[372] = 0;
 buffer[373] = 0;
 buffer[374] = 0;
 buffer[375] = 0;
 buffer[376] = 0;
 buffer[377] = 0;
 buffer[378] = 0;
 buffer[379] = 0;
 buffer[380] = 0;
 buffer[381] = 0;
 buffer[382] = 0;
 buffer[383] = 0;
 buffer[384] = 0;
 buffer[385] = 0;
 buffer[386] = 0;
 buffer[387] = 0;
 buffer[388] = 0;
 buffer[389] = 0;
 buffer[390] = 0;
 buffer[391] = 0;
 buffer[392] = 0;
 buffer[393] = 0;
 buffer[394] = 0;
 buffer[395] = 0;
 buffer[396] = 0;
 buffer[397] = 0;
 buffer[398] = 0;
 buffer[399] = 0;
 buffer[400] = 0;
 buffer[401] = 0;
 buffer[402] = 0;
 buffer[403] = 0;
 buffer[404] = 0;
 buffer[405] = 0;
 buffer[406] = 0;
 buffer[407] = 0;
 buffer[408] = 0;
 buffer[409] = 0;
 buffer[410] = 0;
 buffer[411] = 0;
 buffer[412] = 0;
 buffer[413] = 0;
 buffer[414] = 0;
 buffer[415] = 0;
 buffer[416] = 0;
 buffer[417] = 0;
 buffer[418] = 0;
 buffer[419] = 0;
 buffer[420] = 0;
 buffer[421] = 0;
 buffer[422] = 0;
 buffer[423] = 0;
 buffer[424] = 0;
 buffer[425] = 0;
 buffer[426] = 0;
 buffer[427] = 0;
 buffer[428] = 0;
 buffer[429] = 0;
 buffer[430] = 0;
 buffer[431] = 0;
 buffer[432] = 0;
 buffer[433] = 0;
 buffer[434] = 0;
 buffer[435] = 0;
 buffer[436] = 0;
 buffer[437] = 0;
 buffer[438] = 0;
 buffer[439] = 0;
 buffer[440] = 0;
 buffer[441] = 0;
 buffer[442] = 0;
 buffer[443] = 0;
 buffer[444] = 0;
 buffer[445] = 0;
 buffer[446] = 0;
 buffer[447] = 0;
 buffer[448] = 0;
 buffer[449] = 0;
 buffer[450] = 0;
 buffer[451] = 0;
 buffer[452] = 0;
 buffer[453] = 0;
 buffer[454] = 0;
 buffer[455] = 0;
 buffer[456] = 0;
 buffer[457] = 0;
 buffer[458] = 0;
 buffer[459] = 0;
 buffer[460] = 0;
 buffer[461] = 0;
 buffer[462] = 0;
 buffer[463] = 0;
 buffer[464] = 0;
 buffer[465] = 0;
 buffer[466] = 0;
 buffer[467] = 0;
 buffer[468] = 0;
 buffer[469] = 0;
 buffer[470] = 0;
 buffer[471] = 0;
 buffer[472] = 0;
 buffer[473] = 0;
 buffer[474] = 0;
 buffer[475] = 0;
 buffer[476] = 0;
 buffer[477] = 0;
 buffer[478] = 0;
 buffer[479] = 0;
 buffer[480] = 0;
 buffer[481] = 0;
 buffer[482] = 0;
 buffer[483] = 0;
 buffer[484] = 0;
 buffer[485] = 0;
 buffer[486] = 0;
 buffer[487] = 0;
 buffer[488] = 0;
 buffer[489] = 0;
 buffer[490] = 0;
 buffer[491] = 0;
 buffer[492] = 0;
 buffer[493] = 0;
 buffer[494] = 0;
 buffer[495] = 0;
 buffer[496] = 0;
 buffer[497] = 0;
 buffer[498] = 0;
 buffer[499] = 0;
 buffer[500] = 0;
 buffer[501] = 0;
 buffer[502] = 0;
 buffer[503] = 0;
 buffer[504] = 0;
 buffer[505] = 0;
 buffer[506] = 0;
 buffer[507] = 0;
 buffer[508] = 0;
 buffer[509] = 0;
 buffer[510] = 0;
 buffer[511] = 0;
end

endmodule

module M_tilemap_mem_tiles(
input      [10:0]                in_tiles_addr0,
output reg  [17:0]     out_tiles_rdata0,
output reg  [17:0]     out_tiles_rdata1,
input      [0:0]             in_tiles_wenable1,
input      [17:0]                 in_tiles_wdata1,
input      [10:0]                in_tiles_addr1,
input      clock0,
input      clock1
);
reg  [17:0] buffer[1343:0];
always @(posedge clock0) begin
  out_tiles_rdata0 <= buffer[in_tiles_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_wenable1) begin
    buffer[in_tiles_addr1] <= in_tiles_wdata1;
  end
end
initial begin
 buffer[0] = 18'b100000000000000000;
 buffer[1] = 18'b100000000000000000;
 buffer[2] = 18'b100000000000000000;
 buffer[3] = 18'b100000000000000000;
 buffer[4] = 18'b100000000000000000;
 buffer[5] = 18'b100000000000000000;
 buffer[6] = 18'b100000000000000000;
 buffer[7] = 18'b100000000000000000;
 buffer[8] = 18'b100000000000000000;
 buffer[9] = 18'b100000000000000000;
 buffer[10] = 18'b100000000000000000;
 buffer[11] = 18'b100000000000000000;
 buffer[12] = 18'b100000000000000000;
 buffer[13] = 18'b100000000000000000;
 buffer[14] = 18'b100000000000000000;
 buffer[15] = 18'b100000000000000000;
 buffer[16] = 18'b100000000000000000;
 buffer[17] = 18'b100000000000000000;
 buffer[18] = 18'b100000000000000000;
 buffer[19] = 18'b100000000000000000;
 buffer[20] = 18'b100000000000000000;
 buffer[21] = 18'b100000000000000000;
 buffer[22] = 18'b100000000000000000;
 buffer[23] = 18'b100000000000000000;
 buffer[24] = 18'b100000000000000000;
 buffer[25] = 18'b100000000000000000;
 buffer[26] = 18'b100000000000000000;
 buffer[27] = 18'b100000000000000000;
 buffer[28] = 18'b100000000000000000;
 buffer[29] = 18'b100000000000000000;
 buffer[30] = 18'b100000000000000000;
 buffer[31] = 18'b100000000000000000;
 buffer[32] = 18'b100000000000000000;
 buffer[33] = 18'b100000000000000000;
 buffer[34] = 18'b100000000000000000;
 buffer[35] = 18'b100000000000000000;
 buffer[36] = 18'b100000000000000000;
 buffer[37] = 18'b100000000000000000;
 buffer[38] = 18'b100000000000000000;
 buffer[39] = 18'b100000000000000000;
 buffer[40] = 18'b100000000000000000;
 buffer[41] = 18'b100000000000000000;
 buffer[42] = 18'b100000000000000000;
 buffer[43] = 18'b100000000000000000;
 buffer[44] = 18'b100000000000000000;
 buffer[45] = 18'b100000000000000000;
 buffer[46] = 18'b100000000000000000;
 buffer[47] = 18'b100000000000000000;
 buffer[48] = 18'b100000000000000000;
 buffer[49] = 18'b100000000000000000;
 buffer[50] = 18'b100000000000000000;
 buffer[51] = 18'b100000000000000000;
 buffer[52] = 18'b100000000000000000;
 buffer[53] = 18'b100000000000000000;
 buffer[54] = 18'b100000000000000000;
 buffer[55] = 18'b100000000000000000;
 buffer[56] = 18'b100000000000000000;
 buffer[57] = 18'b100000000000000000;
 buffer[58] = 18'b100000000000000000;
 buffer[59] = 18'b100000000000000000;
 buffer[60] = 18'b100000000000000000;
 buffer[61] = 18'b100000000000000000;
 buffer[62] = 18'b100000000000000000;
 buffer[63] = 18'b100000000000000000;
 buffer[64] = 18'b100000000000000000;
 buffer[65] = 18'b100000000000000000;
 buffer[66] = 18'b100000000000000000;
 buffer[67] = 18'b100000000000000000;
 buffer[68] = 18'b100000000000000000;
 buffer[69] = 18'b100000000000000000;
 buffer[70] = 18'b100000000000000000;
 buffer[71] = 18'b100000000000000000;
 buffer[72] = 18'b100000000000000000;
 buffer[73] = 18'b100000000000000000;
 buffer[74] = 18'b100000000000000000;
 buffer[75] = 18'b100000000000000000;
 buffer[76] = 18'b100000000000000000;
 buffer[77] = 18'b100000000000000000;
 buffer[78] = 18'b100000000000000000;
 buffer[79] = 18'b100000000000000000;
 buffer[80] = 18'b100000000000000000;
 buffer[81] = 18'b100000000000000000;
 buffer[82] = 18'b100000000000000000;
 buffer[83] = 18'b100000000000000000;
 buffer[84] = 18'b100000000000000000;
 buffer[85] = 18'b100000000000000000;
 buffer[86] = 18'b100000000000000000;
 buffer[87] = 18'b100000000000000000;
 buffer[88] = 18'b100000000000000000;
 buffer[89] = 18'b100000000000000000;
 buffer[90] = 18'b100000000000000000;
 buffer[91] = 18'b100000000000000000;
 buffer[92] = 18'b100000000000000000;
 buffer[93] = 18'b100000000000000000;
 buffer[94] = 18'b100000000000000000;
 buffer[95] = 18'b100000000000000000;
 buffer[96] = 18'b100000000000000000;
 buffer[97] = 18'b100000000000000000;
 buffer[98] = 18'b100000000000000000;
 buffer[99] = 18'b100000000000000000;
 buffer[100] = 18'b100000000000000000;
 buffer[101] = 18'b100000000000000000;
 buffer[102] = 18'b100000000000000000;
 buffer[103] = 18'b100000000000000000;
 buffer[104] = 18'b100000000000000000;
 buffer[105] = 18'b100000000000000000;
 buffer[106] = 18'b100000000000000000;
 buffer[107] = 18'b100000000000000000;
 buffer[108] = 18'b100000000000000000;
 buffer[109] = 18'b100000000000000000;
 buffer[110] = 18'b100000000000000000;
 buffer[111] = 18'b100000000000000000;
 buffer[112] = 18'b100000000000000000;
 buffer[113] = 18'b100000000000000000;
 buffer[114] = 18'b100000000000000000;
 buffer[115] = 18'b100000000000000000;
 buffer[116] = 18'b100000000000000000;
 buffer[117] = 18'b100000000000000000;
 buffer[118] = 18'b100000000000000000;
 buffer[119] = 18'b100000000000000000;
 buffer[120] = 18'b100000000000000000;
 buffer[121] = 18'b100000000000000000;
 buffer[122] = 18'b100000000000000000;
 buffer[123] = 18'b100000000000000000;
 buffer[124] = 18'b100000000000000000;
 buffer[125] = 18'b100000000000000000;
 buffer[126] = 18'b100000000000000000;
 buffer[127] = 18'b100000000000000000;
 buffer[128] = 18'b100000000000000000;
 buffer[129] = 18'b100000000000000000;
 buffer[130] = 18'b100000000000000000;
 buffer[131] = 18'b100000000000000000;
 buffer[132] = 18'b100000000000000000;
 buffer[133] = 18'b100000000000000000;
 buffer[134] = 18'b100000000000000000;
 buffer[135] = 18'b100000000000000000;
 buffer[136] = 18'b100000000000000000;
 buffer[137] = 18'b100000000000000000;
 buffer[138] = 18'b100000000000000000;
 buffer[139] = 18'b100000000000000000;
 buffer[140] = 18'b100000000000000000;
 buffer[141] = 18'b100000000000000000;
 buffer[142] = 18'b100000000000000000;
 buffer[143] = 18'b100000000000000000;
 buffer[144] = 18'b100000000000000000;
 buffer[145] = 18'b100000000000000000;
 buffer[146] = 18'b100000000000000000;
 buffer[147] = 18'b100000000000000000;
 buffer[148] = 18'b100000000000000000;
 buffer[149] = 18'b100000000000000000;
 buffer[150] = 18'b100000000000000000;
 buffer[151] = 18'b100000000000000000;
 buffer[152] = 18'b100000000000000000;
 buffer[153] = 18'b100000000000000000;
 buffer[154] = 18'b100000000000000000;
 buffer[155] = 18'b100000000000000000;
 buffer[156] = 18'b100000000000000000;
 buffer[157] = 18'b100000000000000000;
 buffer[158] = 18'b100000000000000000;
 buffer[159] = 18'b100000000000000000;
 buffer[160] = 18'b100000000000000000;
 buffer[161] = 18'b100000000000000000;
 buffer[162] = 18'b100000000000000000;
 buffer[163] = 18'b100000000000000000;
 buffer[164] = 18'b100000000000000000;
 buffer[165] = 18'b100000000000000000;
 buffer[166] = 18'b100000000000000000;
 buffer[167] = 18'b100000000000000000;
 buffer[168] = 18'b100000000000000000;
 buffer[169] = 18'b100000000000000000;
 buffer[170] = 18'b100000000000000000;
 buffer[171] = 18'b100000000000000000;
 buffer[172] = 18'b100000000000000000;
 buffer[173] = 18'b100000000000000000;
 buffer[174] = 18'b100000000000000000;
 buffer[175] = 18'b100000000000000000;
 buffer[176] = 18'b100000000000000000;
 buffer[177] = 18'b100000000000000000;
 buffer[178] = 18'b100000000000000000;
 buffer[179] = 18'b100000000000000000;
 buffer[180] = 18'b100000000000000000;
 buffer[181] = 18'b100000000000000000;
 buffer[182] = 18'b100000000000000000;
 buffer[183] = 18'b100000000000000000;
 buffer[184] = 18'b100000000000000000;
 buffer[185] = 18'b100000000000000000;
 buffer[186] = 18'b100000000000000000;
 buffer[187] = 18'b100000000000000000;
 buffer[188] = 18'b100000000000000000;
 buffer[189] = 18'b100000000000000000;
 buffer[190] = 18'b100000000000000000;
 buffer[191] = 18'b100000000000000000;
 buffer[192] = 18'b100000000000000000;
 buffer[193] = 18'b100000000000000000;
 buffer[194] = 18'b100000000000000000;
 buffer[195] = 18'b100000000000000000;
 buffer[196] = 18'b100000000000000000;
 buffer[197] = 18'b100000000000000000;
 buffer[198] = 18'b100000000000000000;
 buffer[199] = 18'b100000000000000000;
 buffer[200] = 18'b100000000000000000;
 buffer[201] = 18'b100000000000000000;
 buffer[202] = 18'b100000000000000000;
 buffer[203] = 18'b100000000000000000;
 buffer[204] = 18'b100000000000000000;
 buffer[205] = 18'b100000000000000000;
 buffer[206] = 18'b100000000000000000;
 buffer[207] = 18'b100000000000000000;
 buffer[208] = 18'b100000000000000000;
 buffer[209] = 18'b100000000000000000;
 buffer[210] = 18'b100000000000000000;
 buffer[211] = 18'b100000000000000000;
 buffer[212] = 18'b100000000000000000;
 buffer[213] = 18'b100000000000000000;
 buffer[214] = 18'b100000000000000000;
 buffer[215] = 18'b100000000000000000;
 buffer[216] = 18'b100000000000000000;
 buffer[217] = 18'b100000000000000000;
 buffer[218] = 18'b100000000000000000;
 buffer[219] = 18'b100000000000000000;
 buffer[220] = 18'b100000000000000000;
 buffer[221] = 18'b100000000000000000;
 buffer[222] = 18'b100000000000000000;
 buffer[223] = 18'b100000000000000000;
 buffer[224] = 18'b100000000000000000;
 buffer[225] = 18'b100000000000000000;
 buffer[226] = 18'b100000000000000000;
 buffer[227] = 18'b100000000000000000;
 buffer[228] = 18'b100000000000000000;
 buffer[229] = 18'b100000000000000000;
 buffer[230] = 18'b100000000000000000;
 buffer[231] = 18'b100000000000000000;
 buffer[232] = 18'b100000000000000000;
 buffer[233] = 18'b100000000000000000;
 buffer[234] = 18'b100000000000000000;
 buffer[235] = 18'b100000000000000000;
 buffer[236] = 18'b100000000000000000;
 buffer[237] = 18'b100000000000000000;
 buffer[238] = 18'b100000000000000000;
 buffer[239] = 18'b100000000000000000;
 buffer[240] = 18'b100000000000000000;
 buffer[241] = 18'b100000000000000000;
 buffer[242] = 18'b100000000000000000;
 buffer[243] = 18'b100000000000000000;
 buffer[244] = 18'b100000000000000000;
 buffer[245] = 18'b100000000000000000;
 buffer[246] = 18'b100000000000000000;
 buffer[247] = 18'b100000000000000000;
 buffer[248] = 18'b100000000000000000;
 buffer[249] = 18'b100000000000000000;
 buffer[250] = 18'b100000000000000000;
 buffer[251] = 18'b100000000000000000;
 buffer[252] = 18'b100000000000000000;
 buffer[253] = 18'b100000000000000000;
 buffer[254] = 18'b100000000000000000;
 buffer[255] = 18'b100000000000000000;
 buffer[256] = 18'b100000000000000000;
 buffer[257] = 18'b100000000000000000;
 buffer[258] = 18'b100000000000000000;
 buffer[259] = 18'b100000000000000000;
 buffer[260] = 18'b100000000000000000;
 buffer[261] = 18'b100000000000000000;
 buffer[262] = 18'b100000000000000000;
 buffer[263] = 18'b100000000000000000;
 buffer[264] = 18'b100000000000000000;
 buffer[265] = 18'b100000000000000000;
 buffer[266] = 18'b100000000000000000;
 buffer[267] = 18'b100000000000000000;
 buffer[268] = 18'b100000000000000000;
 buffer[269] = 18'b100000000000000000;
 buffer[270] = 18'b100000000000000000;
 buffer[271] = 18'b100000000000000000;
 buffer[272] = 18'b100000000000000000;
 buffer[273] = 18'b100000000000000000;
 buffer[274] = 18'b100000000000000000;
 buffer[275] = 18'b100000000000000000;
 buffer[276] = 18'b100000000000000000;
 buffer[277] = 18'b100000000000000000;
 buffer[278] = 18'b100000000000000000;
 buffer[279] = 18'b100000000000000000;
 buffer[280] = 18'b100000000000000000;
 buffer[281] = 18'b100000000000000000;
 buffer[282] = 18'b100000000000000000;
 buffer[283] = 18'b100000000000000000;
 buffer[284] = 18'b100000000000000000;
 buffer[285] = 18'b100000000000000000;
 buffer[286] = 18'b100000000000000000;
 buffer[287] = 18'b100000000000000000;
 buffer[288] = 18'b100000000000000000;
 buffer[289] = 18'b100000000000000000;
 buffer[290] = 18'b100000000000000000;
 buffer[291] = 18'b100000000000000000;
 buffer[292] = 18'b100000000000000000;
 buffer[293] = 18'b100000000000000000;
 buffer[294] = 18'b100000000000000000;
 buffer[295] = 18'b100000000000000000;
 buffer[296] = 18'b100000000000000000;
 buffer[297] = 18'b100000000000000000;
 buffer[298] = 18'b100000000000000000;
 buffer[299] = 18'b100000000000000000;
 buffer[300] = 18'b100000000000000000;
 buffer[301] = 18'b100000000000000000;
 buffer[302] = 18'b100000000000000000;
 buffer[303] = 18'b100000000000000000;
 buffer[304] = 18'b100000000000000000;
 buffer[305] = 18'b100000000000000000;
 buffer[306] = 18'b100000000000000000;
 buffer[307] = 18'b100000000000000000;
 buffer[308] = 18'b100000000000000000;
 buffer[309] = 18'b100000000000000000;
 buffer[310] = 18'b100000000000000000;
 buffer[311] = 18'b100000000000000000;
 buffer[312] = 18'b100000000000000000;
 buffer[313] = 18'b100000000000000000;
 buffer[314] = 18'b100000000000000000;
 buffer[315] = 18'b100000000000000000;
 buffer[316] = 18'b100000000000000000;
 buffer[317] = 18'b100000000000000000;
 buffer[318] = 18'b100000000000000000;
 buffer[319] = 18'b100000000000000000;
 buffer[320] = 18'b100000000000000000;
 buffer[321] = 18'b100000000000000000;
 buffer[322] = 18'b100000000000000000;
 buffer[323] = 18'b100000000000000000;
 buffer[324] = 18'b100000000000000000;
 buffer[325] = 18'b100000000000000000;
 buffer[326] = 18'b100000000000000000;
 buffer[327] = 18'b100000000000000000;
 buffer[328] = 18'b100000000000000000;
 buffer[329] = 18'b100000000000000000;
 buffer[330] = 18'b100000000000000000;
 buffer[331] = 18'b100000000000000000;
 buffer[332] = 18'b100000000000000000;
 buffer[333] = 18'b100000000000000000;
 buffer[334] = 18'b100000000000000000;
 buffer[335] = 18'b100000000000000000;
 buffer[336] = 18'b100000000000000000;
 buffer[337] = 18'b100000000000000000;
 buffer[338] = 18'b100000000000000000;
 buffer[339] = 18'b100000000000000000;
 buffer[340] = 18'b100000000000000000;
 buffer[341] = 18'b100000000000000000;
 buffer[342] = 18'b100000000000000000;
 buffer[343] = 18'b100000000000000000;
 buffer[344] = 18'b100000000000000000;
 buffer[345] = 18'b100000000000000000;
 buffer[346] = 18'b100000000000000000;
 buffer[347] = 18'b100000000000000000;
 buffer[348] = 18'b100000000000000000;
 buffer[349] = 18'b100000000000000000;
 buffer[350] = 18'b100000000000000000;
 buffer[351] = 18'b100000000000000000;
 buffer[352] = 18'b100000000000000000;
 buffer[353] = 18'b100000000000000000;
 buffer[354] = 18'b100000000000000000;
 buffer[355] = 18'b100000000000000000;
 buffer[356] = 18'b100000000000000000;
 buffer[357] = 18'b100000000000000000;
 buffer[358] = 18'b100000000000000000;
 buffer[359] = 18'b100000000000000000;
 buffer[360] = 18'b100000000000000000;
 buffer[361] = 18'b100000000000000000;
 buffer[362] = 18'b100000000000000000;
 buffer[363] = 18'b100000000000000000;
 buffer[364] = 18'b100000000000000000;
 buffer[365] = 18'b100000000000000000;
 buffer[366] = 18'b100000000000000000;
 buffer[367] = 18'b100000000000000000;
 buffer[368] = 18'b100000000000000000;
 buffer[369] = 18'b100000000000000000;
 buffer[370] = 18'b100000000000000000;
 buffer[371] = 18'b100000000000000000;
 buffer[372] = 18'b100000000000000000;
 buffer[373] = 18'b100000000000000000;
 buffer[374] = 18'b100000000000000000;
 buffer[375] = 18'b100000000000000000;
 buffer[376] = 18'b100000000000000000;
 buffer[377] = 18'b100000000000000000;
 buffer[378] = 18'b100000000000000000;
 buffer[379] = 18'b100000000000000000;
 buffer[380] = 18'b100000000000000000;
 buffer[381] = 18'b100000000000000000;
 buffer[382] = 18'b100000000000000000;
 buffer[383] = 18'b100000000000000000;
 buffer[384] = 18'b100000000000000000;
 buffer[385] = 18'b100000000000000000;
 buffer[386] = 18'b100000000000000000;
 buffer[387] = 18'b100000000000000000;
 buffer[388] = 18'b100000000000000000;
 buffer[389] = 18'b100000000000000000;
 buffer[390] = 18'b100000000000000000;
 buffer[391] = 18'b100000000000000000;
 buffer[392] = 18'b100000000000000000;
 buffer[393] = 18'b100000000000000000;
 buffer[394] = 18'b100000000000000000;
 buffer[395] = 18'b100000000000000000;
 buffer[396] = 18'b100000000000000000;
 buffer[397] = 18'b100000000000000000;
 buffer[398] = 18'b100000000000000000;
 buffer[399] = 18'b100000000000000000;
 buffer[400] = 18'b100000000000000000;
 buffer[401] = 18'b100000000000000000;
 buffer[402] = 18'b100000000000000000;
 buffer[403] = 18'b100000000000000000;
 buffer[404] = 18'b100000000000000000;
 buffer[405] = 18'b100000000000000000;
 buffer[406] = 18'b100000000000000000;
 buffer[407] = 18'b100000000000000000;
 buffer[408] = 18'b100000000000000000;
 buffer[409] = 18'b100000000000000000;
 buffer[410] = 18'b100000000000000000;
 buffer[411] = 18'b100000000000000000;
 buffer[412] = 18'b100000000000000000;
 buffer[413] = 18'b100000000000000000;
 buffer[414] = 18'b100000000000000000;
 buffer[415] = 18'b100000000000000000;
 buffer[416] = 18'b100000000000000000;
 buffer[417] = 18'b100000000000000000;
 buffer[418] = 18'b100000000000000000;
 buffer[419] = 18'b100000000000000000;
 buffer[420] = 18'b100000000000000000;
 buffer[421] = 18'b100000000000000000;
 buffer[422] = 18'b100000000000000000;
 buffer[423] = 18'b100000000000000000;
 buffer[424] = 18'b100000000000000000;
 buffer[425] = 18'b100000000000000000;
 buffer[426] = 18'b100000000000000000;
 buffer[427] = 18'b100000000000000000;
 buffer[428] = 18'b100000000000000000;
 buffer[429] = 18'b100000000000000000;
 buffer[430] = 18'b100000000000000000;
 buffer[431] = 18'b100000000000000000;
 buffer[432] = 18'b100000000000000000;
 buffer[433] = 18'b100000000000000000;
 buffer[434] = 18'b100000000000000000;
 buffer[435] = 18'b100000000000000000;
 buffer[436] = 18'b100000000000000000;
 buffer[437] = 18'b100000000000000000;
 buffer[438] = 18'b100000000000000000;
 buffer[439] = 18'b100000000000000000;
 buffer[440] = 18'b100000000000000000;
 buffer[441] = 18'b100000000000000000;
 buffer[442] = 18'b100000000000000000;
 buffer[443] = 18'b100000000000000000;
 buffer[444] = 18'b100000000000000000;
 buffer[445] = 18'b100000000000000000;
 buffer[446] = 18'b100000000000000000;
 buffer[447] = 18'b100000000000000000;
 buffer[448] = 18'b100000000000000000;
 buffer[449] = 18'b100000000000000000;
 buffer[450] = 18'b100000000000000000;
 buffer[451] = 18'b100000000000000000;
 buffer[452] = 18'b100000000000000000;
 buffer[453] = 18'b100000000000000000;
 buffer[454] = 18'b100000000000000000;
 buffer[455] = 18'b100000000000000000;
 buffer[456] = 18'b100000000000000000;
 buffer[457] = 18'b100000000000000000;
 buffer[458] = 18'b100000000000000000;
 buffer[459] = 18'b100000000000000000;
 buffer[460] = 18'b100000000000000000;
 buffer[461] = 18'b100000000000000000;
 buffer[462] = 18'b100000000000000000;
 buffer[463] = 18'b100000000000000000;
 buffer[464] = 18'b100000000000000000;
 buffer[465] = 18'b100000000000000000;
 buffer[466] = 18'b100000000000000000;
 buffer[467] = 18'b100000000000000000;
 buffer[468] = 18'b100000000000000000;
 buffer[469] = 18'b100000000000000000;
 buffer[470] = 18'b100000000000000000;
 buffer[471] = 18'b100000000000000000;
 buffer[472] = 18'b100000000000000000;
 buffer[473] = 18'b100000000000000000;
 buffer[474] = 18'b100000000000000000;
 buffer[475] = 18'b100000000000000000;
 buffer[476] = 18'b100000000000000000;
 buffer[477] = 18'b100000000000000000;
 buffer[478] = 18'b100000000000000000;
 buffer[479] = 18'b100000000000000000;
 buffer[480] = 18'b100000000000000000;
 buffer[481] = 18'b100000000000000000;
 buffer[482] = 18'b100000000000000000;
 buffer[483] = 18'b100000000000000000;
 buffer[484] = 18'b100000000000000000;
 buffer[485] = 18'b100000000000000000;
 buffer[486] = 18'b100000000000000000;
 buffer[487] = 18'b100000000000000000;
 buffer[488] = 18'b100000000000000000;
 buffer[489] = 18'b100000000000000000;
 buffer[490] = 18'b100000000000000000;
 buffer[491] = 18'b100000000000000000;
 buffer[492] = 18'b100000000000000000;
 buffer[493] = 18'b100000000000000000;
 buffer[494] = 18'b100000000000000000;
 buffer[495] = 18'b100000000000000000;
 buffer[496] = 18'b100000000000000000;
 buffer[497] = 18'b100000000000000000;
 buffer[498] = 18'b100000000000000000;
 buffer[499] = 18'b100000000000000000;
 buffer[500] = 18'b100000000000000000;
 buffer[501] = 18'b100000000000000000;
 buffer[502] = 18'b100000000000000000;
 buffer[503] = 18'b100000000000000000;
 buffer[504] = 18'b100000000000000000;
 buffer[505] = 18'b100000000000000000;
 buffer[506] = 18'b100000000000000000;
 buffer[507] = 18'b100000000000000000;
 buffer[508] = 18'b100000000000000000;
 buffer[509] = 18'b100000000000000000;
 buffer[510] = 18'b100000000000000000;
 buffer[511] = 18'b100000000000000000;
 buffer[512] = 18'b100000000000000000;
 buffer[513] = 18'b100000000000000000;
 buffer[514] = 18'b100000000000000000;
 buffer[515] = 18'b100000000000000000;
 buffer[516] = 18'b100000000000000000;
 buffer[517] = 18'b100000000000000000;
 buffer[518] = 18'b100000000000000000;
 buffer[519] = 18'b100000000000000000;
 buffer[520] = 18'b100000000000000000;
 buffer[521] = 18'b100000000000000000;
 buffer[522] = 18'b100000000000000000;
 buffer[523] = 18'b100000000000000000;
 buffer[524] = 18'b100000000000000000;
 buffer[525] = 18'b100000000000000000;
 buffer[526] = 18'b100000000000000000;
 buffer[527] = 18'b100000000000000000;
 buffer[528] = 18'b100000000000000000;
 buffer[529] = 18'b100000000000000000;
 buffer[530] = 18'b100000000000000000;
 buffer[531] = 18'b100000000000000000;
 buffer[532] = 18'b100000000000000000;
 buffer[533] = 18'b100000000000000000;
 buffer[534] = 18'b100000000000000000;
 buffer[535] = 18'b100000000000000000;
 buffer[536] = 18'b100000000000000000;
 buffer[537] = 18'b100000000000000000;
 buffer[538] = 18'b100000000000000000;
 buffer[539] = 18'b100000000000000000;
 buffer[540] = 18'b100000000000000000;
 buffer[541] = 18'b100000000000000000;
 buffer[542] = 18'b100000000000000000;
 buffer[543] = 18'b100000000000000000;
 buffer[544] = 18'b100000000000000000;
 buffer[545] = 18'b100000000000000000;
 buffer[546] = 18'b100000000000000000;
 buffer[547] = 18'b100000000000000000;
 buffer[548] = 18'b100000000000000000;
 buffer[549] = 18'b100000000000000000;
 buffer[550] = 18'b100000000000000000;
 buffer[551] = 18'b100000000000000000;
 buffer[552] = 18'b100000000000000000;
 buffer[553] = 18'b100000000000000000;
 buffer[554] = 18'b100000000000000000;
 buffer[555] = 18'b100000000000000000;
 buffer[556] = 18'b100000000000000000;
 buffer[557] = 18'b100000000000000000;
 buffer[558] = 18'b100000000000000000;
 buffer[559] = 18'b100000000000000000;
 buffer[560] = 18'b100000000000000000;
 buffer[561] = 18'b100000000000000000;
 buffer[562] = 18'b100000000000000000;
 buffer[563] = 18'b100000000000000000;
 buffer[564] = 18'b100000000000000000;
 buffer[565] = 18'b100000000000000000;
 buffer[566] = 18'b100000000000000000;
 buffer[567] = 18'b100000000000000000;
 buffer[568] = 18'b100000000000000000;
 buffer[569] = 18'b100000000000000000;
 buffer[570] = 18'b100000000000000000;
 buffer[571] = 18'b100000000000000000;
 buffer[572] = 18'b100000000000000000;
 buffer[573] = 18'b100000000000000000;
 buffer[574] = 18'b100000000000000000;
 buffer[575] = 18'b100000000000000000;
 buffer[576] = 18'b100000000000000000;
 buffer[577] = 18'b100000000000000000;
 buffer[578] = 18'b100000000000000000;
 buffer[579] = 18'b100000000000000000;
 buffer[580] = 18'b100000000000000000;
 buffer[581] = 18'b100000000000000000;
 buffer[582] = 18'b100000000000000000;
 buffer[583] = 18'b100000000000000000;
 buffer[584] = 18'b100000000000000000;
 buffer[585] = 18'b100000000000000000;
 buffer[586] = 18'b100000000000000000;
 buffer[587] = 18'b100000000000000000;
 buffer[588] = 18'b100000000000000000;
 buffer[589] = 18'b100000000000000000;
 buffer[590] = 18'b100000000000000000;
 buffer[591] = 18'b100000000000000000;
 buffer[592] = 18'b100000000000000000;
 buffer[593] = 18'b100000000000000000;
 buffer[594] = 18'b100000000000000000;
 buffer[595] = 18'b100000000000000000;
 buffer[596] = 18'b100000000000000000;
 buffer[597] = 18'b100000000000000000;
 buffer[598] = 18'b100000000000000000;
 buffer[599] = 18'b100000000000000000;
 buffer[600] = 18'b100000000000000000;
 buffer[601] = 18'b100000000000000000;
 buffer[602] = 18'b100000000000000000;
 buffer[603] = 18'b100000000000000000;
 buffer[604] = 18'b100000000000000000;
 buffer[605] = 18'b100000000000000000;
 buffer[606] = 18'b100000000000000000;
 buffer[607] = 18'b100000000000000000;
 buffer[608] = 18'b100000000000000000;
 buffer[609] = 18'b100000000000000000;
 buffer[610] = 18'b100000000000000000;
 buffer[611] = 18'b100000000000000000;
 buffer[612] = 18'b100000000000000000;
 buffer[613] = 18'b100000000000000000;
 buffer[614] = 18'b100000000000000000;
 buffer[615] = 18'b100000000000000000;
 buffer[616] = 18'b100000000000000000;
 buffer[617] = 18'b100000000000000000;
 buffer[618] = 18'b100000000000000000;
 buffer[619] = 18'b100000000000000000;
 buffer[620] = 18'b100000000000000000;
 buffer[621] = 18'b100000000000000000;
 buffer[622] = 18'b100000000000000000;
 buffer[623] = 18'b100000000000000000;
 buffer[624] = 18'b100000000000000000;
 buffer[625] = 18'b100000000000000000;
 buffer[626] = 18'b100000000000000000;
 buffer[627] = 18'b100000000000000000;
 buffer[628] = 18'b100000000000000000;
 buffer[629] = 18'b100000000000000000;
 buffer[630] = 18'b100000000000000000;
 buffer[631] = 18'b100000000000000000;
 buffer[632] = 18'b100000000000000000;
 buffer[633] = 18'b100000000000000000;
 buffer[634] = 18'b100000000000000000;
 buffer[635] = 18'b100000000000000000;
 buffer[636] = 18'b100000000000000000;
 buffer[637] = 18'b100000000000000000;
 buffer[638] = 18'b100000000000000000;
 buffer[639] = 18'b100000000000000000;
 buffer[640] = 18'b100000000000000000;
 buffer[641] = 18'b100000000000000000;
 buffer[642] = 18'b100000000000000000;
 buffer[643] = 18'b100000000000000000;
 buffer[644] = 18'b100000000000000000;
 buffer[645] = 18'b100000000000000000;
 buffer[646] = 18'b100000000000000000;
 buffer[647] = 18'b100000000000000000;
 buffer[648] = 18'b100000000000000000;
 buffer[649] = 18'b100000000000000000;
 buffer[650] = 18'b100000000000000000;
 buffer[651] = 18'b100000000000000000;
 buffer[652] = 18'b100000000000000000;
 buffer[653] = 18'b100000000000000000;
 buffer[654] = 18'b100000000000000000;
 buffer[655] = 18'b100000000000000000;
 buffer[656] = 18'b100000000000000000;
 buffer[657] = 18'b100000000000000000;
 buffer[658] = 18'b100000000000000000;
 buffer[659] = 18'b100000000000000000;
 buffer[660] = 18'b100000000000000000;
 buffer[661] = 18'b100000000000000000;
 buffer[662] = 18'b100000000000000000;
 buffer[663] = 18'b100000000000000000;
 buffer[664] = 18'b100000000000000000;
 buffer[665] = 18'b100000000000000000;
 buffer[666] = 18'b100000000000000000;
 buffer[667] = 18'b100000000000000000;
 buffer[668] = 18'b100000000000000000;
 buffer[669] = 18'b100000000000000000;
 buffer[670] = 18'b100000000000000000;
 buffer[671] = 18'b100000000000000000;
 buffer[672] = 18'b100000000000000000;
 buffer[673] = 18'b100000000000000000;
 buffer[674] = 18'b100000000000000000;
 buffer[675] = 18'b100000000000000000;
 buffer[676] = 18'b100000000000000000;
 buffer[677] = 18'b100000000000000000;
 buffer[678] = 18'b100000000000000000;
 buffer[679] = 18'b100000000000000000;
 buffer[680] = 18'b100000000000000000;
 buffer[681] = 18'b100000000000000000;
 buffer[682] = 18'b100000000000000000;
 buffer[683] = 18'b100000000000000000;
 buffer[684] = 18'b100000000000000000;
 buffer[685] = 18'b100000000000000000;
 buffer[686] = 18'b100000000000000000;
 buffer[687] = 18'b100000000000000000;
 buffer[688] = 18'b100000000000000000;
 buffer[689] = 18'b100000000000000000;
 buffer[690] = 18'b100000000000000000;
 buffer[691] = 18'b100000000000000000;
 buffer[692] = 18'b100000000000000000;
 buffer[693] = 18'b100000000000000000;
 buffer[694] = 18'b100000000000000000;
 buffer[695] = 18'b100000000000000000;
 buffer[696] = 18'b100000000000000000;
 buffer[697] = 18'b100000000000000000;
 buffer[698] = 18'b100000000000000000;
 buffer[699] = 18'b100000000000000000;
 buffer[700] = 18'b100000000000000000;
 buffer[701] = 18'b100000000000000000;
 buffer[702] = 18'b100000000000000000;
 buffer[703] = 18'b100000000000000000;
 buffer[704] = 18'b100000000000000000;
 buffer[705] = 18'b100000000000000000;
 buffer[706] = 18'b100000000000000000;
 buffer[707] = 18'b100000000000000000;
 buffer[708] = 18'b100000000000000000;
 buffer[709] = 18'b100000000000000000;
 buffer[710] = 18'b100000000000000000;
 buffer[711] = 18'b100000000000000000;
 buffer[712] = 18'b100000000000000000;
 buffer[713] = 18'b100000000000000000;
 buffer[714] = 18'b100000000000000000;
 buffer[715] = 18'b100000000000000000;
 buffer[716] = 18'b100000000000000000;
 buffer[717] = 18'b100000000000000000;
 buffer[718] = 18'b100000000000000000;
 buffer[719] = 18'b100000000000000000;
 buffer[720] = 18'b100000000000000000;
 buffer[721] = 18'b100000000000000000;
 buffer[722] = 18'b100000000000000000;
 buffer[723] = 18'b100000000000000000;
 buffer[724] = 18'b100000000000000000;
 buffer[725] = 18'b100000000000000000;
 buffer[726] = 18'b100000000000000000;
 buffer[727] = 18'b100000000000000000;
 buffer[728] = 18'b100000000000000000;
 buffer[729] = 18'b100000000000000000;
 buffer[730] = 18'b100000000000000000;
 buffer[731] = 18'b100000000000000000;
 buffer[732] = 18'b100000000000000000;
 buffer[733] = 18'b100000000000000000;
 buffer[734] = 18'b100000000000000000;
 buffer[735] = 18'b100000000000000000;
 buffer[736] = 18'b100000000000000000;
 buffer[737] = 18'b100000000000000000;
 buffer[738] = 18'b100000000000000000;
 buffer[739] = 18'b100000000000000000;
 buffer[740] = 18'b100000000000000000;
 buffer[741] = 18'b100000000000000000;
 buffer[742] = 18'b100000000000000000;
 buffer[743] = 18'b100000000000000000;
 buffer[744] = 18'b100000000000000000;
 buffer[745] = 18'b100000000000000000;
 buffer[746] = 18'b100000000000000000;
 buffer[747] = 18'b100000000000000000;
 buffer[748] = 18'b100000000000000000;
 buffer[749] = 18'b100000000000000000;
 buffer[750] = 18'b100000000000000000;
 buffer[751] = 18'b100000000000000000;
 buffer[752] = 18'b100000000000000000;
 buffer[753] = 18'b100000000000000000;
 buffer[754] = 18'b100000000000000000;
 buffer[755] = 18'b100000000000000000;
 buffer[756] = 18'b100000000000000000;
 buffer[757] = 18'b100000000000000000;
 buffer[758] = 18'b100000000000000000;
 buffer[759] = 18'b100000000000000000;
 buffer[760] = 18'b100000000000000000;
 buffer[761] = 18'b100000000000000000;
 buffer[762] = 18'b100000000000000000;
 buffer[763] = 18'b100000000000000000;
 buffer[764] = 18'b100000000000000000;
 buffer[765] = 18'b100000000000000000;
 buffer[766] = 18'b100000000000000000;
 buffer[767] = 18'b100000000000000000;
 buffer[768] = 18'b100000000000000000;
 buffer[769] = 18'b100000000000000000;
 buffer[770] = 18'b100000000000000000;
 buffer[771] = 18'b100000000000000000;
 buffer[772] = 18'b100000000000000000;
 buffer[773] = 18'b100000000000000000;
 buffer[774] = 18'b100000000000000000;
 buffer[775] = 18'b100000000000000000;
 buffer[776] = 18'b100000000000000000;
 buffer[777] = 18'b100000000000000000;
 buffer[778] = 18'b100000000000000000;
 buffer[779] = 18'b100000000000000000;
 buffer[780] = 18'b100000000000000000;
 buffer[781] = 18'b100000000000000000;
 buffer[782] = 18'b100000000000000000;
 buffer[783] = 18'b100000000000000000;
 buffer[784] = 18'b100000000000000000;
 buffer[785] = 18'b100000000000000000;
 buffer[786] = 18'b100000000000000000;
 buffer[787] = 18'b100000000000000000;
 buffer[788] = 18'b100000000000000000;
 buffer[789] = 18'b100000000000000000;
 buffer[790] = 18'b100000000000000000;
 buffer[791] = 18'b100000000000000000;
 buffer[792] = 18'b100000000000000000;
 buffer[793] = 18'b100000000000000000;
 buffer[794] = 18'b100000000000000000;
 buffer[795] = 18'b100000000000000000;
 buffer[796] = 18'b100000000000000000;
 buffer[797] = 18'b100000000000000000;
 buffer[798] = 18'b100000000000000000;
 buffer[799] = 18'b100000000000000000;
 buffer[800] = 18'b100000000000000000;
 buffer[801] = 18'b100000000000000000;
 buffer[802] = 18'b100000000000000000;
 buffer[803] = 18'b100000000000000000;
 buffer[804] = 18'b100000000000000000;
 buffer[805] = 18'b100000000000000000;
 buffer[806] = 18'b100000000000000000;
 buffer[807] = 18'b100000000000000000;
 buffer[808] = 18'b100000000000000000;
 buffer[809] = 18'b100000000000000000;
 buffer[810] = 18'b100000000000000000;
 buffer[811] = 18'b100000000000000000;
 buffer[812] = 18'b100000000000000000;
 buffer[813] = 18'b100000000000000000;
 buffer[814] = 18'b100000000000000000;
 buffer[815] = 18'b100000000000000000;
 buffer[816] = 18'b100000000000000000;
 buffer[817] = 18'b100000000000000000;
 buffer[818] = 18'b100000000000000000;
 buffer[819] = 18'b100000000000000000;
 buffer[820] = 18'b100000000000000000;
 buffer[821] = 18'b100000000000000000;
 buffer[822] = 18'b100000000000000000;
 buffer[823] = 18'b100000000000000000;
 buffer[824] = 18'b100000000000000000;
 buffer[825] = 18'b100000000000000000;
 buffer[826] = 18'b100000000000000000;
 buffer[827] = 18'b100000000000000000;
 buffer[828] = 18'b100000000000000000;
 buffer[829] = 18'b100000000000000000;
 buffer[830] = 18'b100000000000000000;
 buffer[831] = 18'b100000000000000000;
 buffer[832] = 18'b100000000000000000;
 buffer[833] = 18'b100000000000000000;
 buffer[834] = 18'b100000000000000000;
 buffer[835] = 18'b100000000000000000;
 buffer[836] = 18'b100000000000000000;
 buffer[837] = 18'b100000000000000000;
 buffer[838] = 18'b100000000000000000;
 buffer[839] = 18'b100000000000000000;
 buffer[840] = 18'b100000000000000000;
 buffer[841] = 18'b100000000000000000;
 buffer[842] = 18'b100000000000000000;
 buffer[843] = 18'b100000000000000000;
 buffer[844] = 18'b100000000000000000;
 buffer[845] = 18'b100000000000000000;
 buffer[846] = 18'b100000000000000000;
 buffer[847] = 18'b100000000000000000;
 buffer[848] = 18'b100000000000000000;
 buffer[849] = 18'b100000000000000000;
 buffer[850] = 18'b100000000000000000;
 buffer[851] = 18'b100000000000000000;
 buffer[852] = 18'b100000000000000000;
 buffer[853] = 18'b100000000000000000;
 buffer[854] = 18'b100000000000000000;
 buffer[855] = 18'b100000000000000000;
 buffer[856] = 18'b100000000000000000;
 buffer[857] = 18'b100000000000000000;
 buffer[858] = 18'b100000000000000000;
 buffer[859] = 18'b100000000000000000;
 buffer[860] = 18'b100000000000000000;
 buffer[861] = 18'b100000000000000000;
 buffer[862] = 18'b100000000000000000;
 buffer[863] = 18'b100000000000000000;
 buffer[864] = 18'b100000000000000000;
 buffer[865] = 18'b100000000000000000;
 buffer[866] = 18'b100000000000000000;
 buffer[867] = 18'b100000000000000000;
 buffer[868] = 18'b100000000000000000;
 buffer[869] = 18'b100000000000000000;
 buffer[870] = 18'b100000000000000000;
 buffer[871] = 18'b100000000000000000;
 buffer[872] = 18'b100000000000000000;
 buffer[873] = 18'b100000000000000000;
 buffer[874] = 18'b100000000000000000;
 buffer[875] = 18'b100000000000000000;
 buffer[876] = 18'b100000000000000000;
 buffer[877] = 18'b100000000000000000;
 buffer[878] = 18'b100000000000000000;
 buffer[879] = 18'b100000000000000000;
 buffer[880] = 18'b100000000000000000;
 buffer[881] = 18'b100000000000000000;
 buffer[882] = 18'b100000000000000000;
 buffer[883] = 18'b100000000000000000;
 buffer[884] = 18'b100000000000000000;
 buffer[885] = 18'b100000000000000000;
 buffer[886] = 18'b100000000000000000;
 buffer[887] = 18'b100000000000000000;
 buffer[888] = 18'b100000000000000000;
 buffer[889] = 18'b100000000000000000;
 buffer[890] = 18'b100000000000000000;
 buffer[891] = 18'b100000000000000000;
 buffer[892] = 18'b100000000000000000;
 buffer[893] = 18'b100000000000000000;
 buffer[894] = 18'b100000000000000000;
 buffer[895] = 18'b100000000000000000;
 buffer[896] = 18'b100000000000000000;
 buffer[897] = 18'b100000000000000000;
 buffer[898] = 18'b100000000000000000;
 buffer[899] = 18'b100000000000000000;
 buffer[900] = 18'b100000000000000000;
 buffer[901] = 18'b100000000000000000;
 buffer[902] = 18'b100000000000000000;
 buffer[903] = 18'b100000000000000000;
 buffer[904] = 18'b100000000000000000;
 buffer[905] = 18'b100000000000000000;
 buffer[906] = 18'b100000000000000000;
 buffer[907] = 18'b100000000000000000;
 buffer[908] = 18'b100000000000000000;
 buffer[909] = 18'b100000000000000000;
 buffer[910] = 18'b100000000000000000;
 buffer[911] = 18'b100000000000000000;
 buffer[912] = 18'b100000000000000000;
 buffer[913] = 18'b100000000000000000;
 buffer[914] = 18'b100000000000000000;
 buffer[915] = 18'b100000000000000000;
 buffer[916] = 18'b100000000000000000;
 buffer[917] = 18'b100000000000000000;
 buffer[918] = 18'b100000000000000000;
 buffer[919] = 18'b100000000000000000;
 buffer[920] = 18'b100000000000000000;
 buffer[921] = 18'b100000000000000000;
 buffer[922] = 18'b100000000000000000;
 buffer[923] = 18'b100000000000000000;
 buffer[924] = 18'b100000000000000000;
 buffer[925] = 18'b100000000000000000;
 buffer[926] = 18'b100000000000000000;
 buffer[927] = 18'b100000000000000000;
 buffer[928] = 18'b100000000000000000;
 buffer[929] = 18'b100000000000000000;
 buffer[930] = 18'b100000000000000000;
 buffer[931] = 18'b100000000000000000;
 buffer[932] = 18'b100000000000000000;
 buffer[933] = 18'b100000000000000000;
 buffer[934] = 18'b100000000000000000;
 buffer[935] = 18'b100000000000000000;
 buffer[936] = 18'b100000000000000000;
 buffer[937] = 18'b100000000000000000;
 buffer[938] = 18'b100000000000000000;
 buffer[939] = 18'b100000000000000000;
 buffer[940] = 18'b100000000000000000;
 buffer[941] = 18'b100000000000000000;
 buffer[942] = 18'b100000000000000000;
 buffer[943] = 18'b100000000000000000;
 buffer[944] = 18'b100000000000000000;
 buffer[945] = 18'b100000000000000000;
 buffer[946] = 18'b100000000000000000;
 buffer[947] = 18'b100000000000000000;
 buffer[948] = 18'b100000000000000000;
 buffer[949] = 18'b100000000000000000;
 buffer[950] = 18'b100000000000000000;
 buffer[951] = 18'b100000000000000000;
 buffer[952] = 18'b100000000000000000;
 buffer[953] = 18'b100000000000000000;
 buffer[954] = 18'b100000000000000000;
 buffer[955] = 18'b100000000000000000;
 buffer[956] = 18'b100000000000000000;
 buffer[957] = 18'b100000000000000000;
 buffer[958] = 18'b100000000000000000;
 buffer[959] = 18'b100000000000000000;
 buffer[960] = 18'b100000000000000000;
 buffer[961] = 18'b100000000000000000;
 buffer[962] = 18'b100000000000000000;
 buffer[963] = 18'b100000000000000000;
 buffer[964] = 18'b100000000000000000;
 buffer[965] = 18'b100000000000000000;
 buffer[966] = 18'b100000000000000000;
 buffer[967] = 18'b100000000000000000;
 buffer[968] = 18'b100000000000000000;
 buffer[969] = 18'b100000000000000000;
 buffer[970] = 18'b100000000000000000;
 buffer[971] = 18'b100000000000000000;
 buffer[972] = 18'b100000000000000000;
 buffer[973] = 18'b100000000000000000;
 buffer[974] = 18'b100000000000000000;
 buffer[975] = 18'b100000000000000000;
 buffer[976] = 18'b100000000000000000;
 buffer[977] = 18'b100000000000000000;
 buffer[978] = 18'b100000000000000000;
 buffer[979] = 18'b100000000000000000;
 buffer[980] = 18'b100000000000000000;
 buffer[981] = 18'b100000000000000000;
 buffer[982] = 18'b100000000000000000;
 buffer[983] = 18'b100000000000000000;
 buffer[984] = 18'b100000000000000000;
 buffer[985] = 18'b100000000000000000;
 buffer[986] = 18'b100000000000000000;
 buffer[987] = 18'b100000000000000000;
 buffer[988] = 18'b100000000000000000;
 buffer[989] = 18'b100000000000000000;
 buffer[990] = 18'b100000000000000000;
 buffer[991] = 18'b100000000000000000;
 buffer[992] = 18'b100000000000000000;
 buffer[993] = 18'b100000000000000000;
 buffer[994] = 18'b100000000000000000;
 buffer[995] = 18'b100000000000000000;
 buffer[996] = 18'b100000000000000000;
 buffer[997] = 18'b100000000000000000;
 buffer[998] = 18'b100000000000000000;
 buffer[999] = 18'b100000000000000000;
 buffer[1000] = 18'b100000000000000000;
 buffer[1001] = 18'b100000000000000000;
 buffer[1002] = 18'b100000000000000000;
 buffer[1003] = 18'b100000000000000000;
 buffer[1004] = 18'b100000000000000000;
 buffer[1005] = 18'b100000000000000000;
 buffer[1006] = 18'b100000000000000000;
 buffer[1007] = 18'b100000000000000000;
 buffer[1008] = 18'b100000000000000000;
 buffer[1009] = 18'b100000000000000000;
 buffer[1010] = 18'b100000000000000000;
 buffer[1011] = 18'b100000000000000000;
 buffer[1012] = 18'b100000000000000000;
 buffer[1013] = 18'b100000000000000000;
 buffer[1014] = 18'b100000000000000000;
 buffer[1015] = 18'b100000000000000000;
 buffer[1016] = 18'b100000000000000000;
 buffer[1017] = 18'b100000000000000000;
 buffer[1018] = 18'b100000000000000000;
 buffer[1019] = 18'b100000000000000000;
 buffer[1020] = 18'b100000000000000000;
 buffer[1021] = 18'b100000000000000000;
 buffer[1022] = 18'b100000000000000000;
 buffer[1023] = 18'b100000000000000000;
 buffer[1024] = 18'b100000000000000000;
 buffer[1025] = 18'b100000000000000000;
 buffer[1026] = 18'b100000000000000000;
 buffer[1027] = 18'b100000000000000000;
 buffer[1028] = 18'b100000000000000000;
 buffer[1029] = 18'b100000000000000000;
 buffer[1030] = 18'b100000000000000000;
 buffer[1031] = 18'b100000000000000000;
 buffer[1032] = 18'b100000000000000000;
 buffer[1033] = 18'b100000000000000000;
 buffer[1034] = 18'b100000000000000000;
 buffer[1035] = 18'b100000000000000000;
 buffer[1036] = 18'b100000000000000000;
 buffer[1037] = 18'b100000000000000000;
 buffer[1038] = 18'b100000000000000000;
 buffer[1039] = 18'b100000000000000000;
 buffer[1040] = 18'b100000000000000000;
 buffer[1041] = 18'b100000000000000000;
 buffer[1042] = 18'b100000000000000000;
 buffer[1043] = 18'b100000000000000000;
 buffer[1044] = 18'b100000000000000000;
 buffer[1045] = 18'b100000000000000000;
 buffer[1046] = 18'b100000000000000000;
 buffer[1047] = 18'b100000000000000000;
 buffer[1048] = 18'b100000000000000000;
 buffer[1049] = 18'b100000000000000000;
 buffer[1050] = 18'b100000000000000000;
 buffer[1051] = 18'b100000000000000000;
 buffer[1052] = 18'b100000000000000000;
 buffer[1053] = 18'b100000000000000000;
 buffer[1054] = 18'b100000000000000000;
 buffer[1055] = 18'b100000000000000000;
 buffer[1056] = 18'b100000000000000000;
 buffer[1057] = 18'b100000000000000000;
 buffer[1058] = 18'b100000000000000000;
 buffer[1059] = 18'b100000000000000000;
 buffer[1060] = 18'b100000000000000000;
 buffer[1061] = 18'b100000000000000000;
 buffer[1062] = 18'b100000000000000000;
 buffer[1063] = 18'b100000000000000000;
 buffer[1064] = 18'b100000000000000000;
 buffer[1065] = 18'b100000000000000000;
 buffer[1066] = 18'b100000000000000000;
 buffer[1067] = 18'b100000000000000000;
 buffer[1068] = 18'b100000000000000000;
 buffer[1069] = 18'b100000000000000000;
 buffer[1070] = 18'b100000000000000000;
 buffer[1071] = 18'b100000000000000000;
 buffer[1072] = 18'b100000000000000000;
 buffer[1073] = 18'b100000000000000000;
 buffer[1074] = 18'b100000000000000000;
 buffer[1075] = 18'b100000000000000000;
 buffer[1076] = 18'b100000000000000000;
 buffer[1077] = 18'b100000000000000000;
 buffer[1078] = 18'b100000000000000000;
 buffer[1079] = 18'b100000000000000000;
 buffer[1080] = 18'b100000000000000000;
 buffer[1081] = 18'b100000000000000000;
 buffer[1082] = 18'b100000000000000000;
 buffer[1083] = 18'b100000000000000000;
 buffer[1084] = 18'b100000000000000000;
 buffer[1085] = 18'b100000000000000000;
 buffer[1086] = 18'b100000000000000000;
 buffer[1087] = 18'b100000000000000000;
 buffer[1088] = 18'b100000000000000000;
 buffer[1089] = 18'b100000000000000000;
 buffer[1090] = 18'b100000000000000000;
 buffer[1091] = 18'b100000000000000000;
 buffer[1092] = 18'b100000000000000000;
 buffer[1093] = 18'b100000000000000000;
 buffer[1094] = 18'b100000000000000000;
 buffer[1095] = 18'b100000000000000000;
 buffer[1096] = 18'b100000000000000000;
 buffer[1097] = 18'b100000000000000000;
 buffer[1098] = 18'b100000000000000000;
 buffer[1099] = 18'b100000000000000000;
 buffer[1100] = 18'b100000000000000000;
 buffer[1101] = 18'b100000000000000000;
 buffer[1102] = 18'b100000000000000000;
 buffer[1103] = 18'b100000000000000000;
 buffer[1104] = 18'b100000000000000000;
 buffer[1105] = 18'b100000000000000000;
 buffer[1106] = 18'b100000000000000000;
 buffer[1107] = 18'b100000000000000000;
 buffer[1108] = 18'b100000000000000000;
 buffer[1109] = 18'b100000000000000000;
 buffer[1110] = 18'b100000000000000000;
 buffer[1111] = 18'b100000000000000000;
 buffer[1112] = 18'b100000000000000000;
 buffer[1113] = 18'b100000000000000000;
 buffer[1114] = 18'b100000000000000000;
 buffer[1115] = 18'b100000000000000000;
 buffer[1116] = 18'b100000000000000000;
 buffer[1117] = 18'b100000000000000000;
 buffer[1118] = 18'b100000000000000000;
 buffer[1119] = 18'b100000000000000000;
 buffer[1120] = 18'b100000000000000000;
 buffer[1121] = 18'b100000000000000000;
 buffer[1122] = 18'b100000000000000000;
 buffer[1123] = 18'b100000000000000000;
 buffer[1124] = 18'b100000000000000000;
 buffer[1125] = 18'b100000000000000000;
 buffer[1126] = 18'b100000000000000000;
 buffer[1127] = 18'b100000000000000000;
 buffer[1128] = 18'b100000000000000000;
 buffer[1129] = 18'b100000000000000000;
 buffer[1130] = 18'b100000000000000000;
 buffer[1131] = 18'b100000000000000000;
 buffer[1132] = 18'b100000000000000000;
 buffer[1133] = 18'b100000000000000000;
 buffer[1134] = 18'b100000000000000000;
 buffer[1135] = 18'b100000000000000000;
 buffer[1136] = 18'b100000000000000000;
 buffer[1137] = 18'b100000000000000000;
 buffer[1138] = 18'b100000000000000000;
 buffer[1139] = 18'b100000000000000000;
 buffer[1140] = 18'b100000000000000000;
 buffer[1141] = 18'b100000000000000000;
 buffer[1142] = 18'b100000000000000000;
 buffer[1143] = 18'b100000000000000000;
 buffer[1144] = 18'b100000000000000000;
 buffer[1145] = 18'b100000000000000000;
 buffer[1146] = 18'b100000000000000000;
 buffer[1147] = 18'b100000000000000000;
 buffer[1148] = 18'b100000000000000000;
 buffer[1149] = 18'b100000000000000000;
 buffer[1150] = 18'b100000000000000000;
 buffer[1151] = 18'b100000000000000000;
 buffer[1152] = 18'b100000000000000000;
 buffer[1153] = 18'b100000000000000000;
 buffer[1154] = 18'b100000000000000000;
 buffer[1155] = 18'b100000000000000000;
 buffer[1156] = 18'b100000000000000000;
 buffer[1157] = 18'b100000000000000000;
 buffer[1158] = 18'b100000000000000000;
 buffer[1159] = 18'b100000000000000000;
 buffer[1160] = 18'b100000000000000000;
 buffer[1161] = 18'b100000000000000000;
 buffer[1162] = 18'b100000000000000000;
 buffer[1163] = 18'b100000000000000000;
 buffer[1164] = 18'b100000000000000000;
 buffer[1165] = 18'b100000000000000000;
 buffer[1166] = 18'b100000000000000000;
 buffer[1167] = 18'b100000000000000000;
 buffer[1168] = 18'b100000000000000000;
 buffer[1169] = 18'b100000000000000000;
 buffer[1170] = 18'b100000000000000000;
 buffer[1171] = 18'b100000000000000000;
 buffer[1172] = 18'b100000000000000000;
 buffer[1173] = 18'b100000000000000000;
 buffer[1174] = 18'b100000000000000000;
 buffer[1175] = 18'b100000000000000000;
 buffer[1176] = 18'b100000000000000000;
 buffer[1177] = 18'b100000000000000000;
 buffer[1178] = 18'b100000000000000000;
 buffer[1179] = 18'b100000000000000000;
 buffer[1180] = 18'b100000000000000000;
 buffer[1181] = 18'b100000000000000000;
 buffer[1182] = 18'b100000000000000000;
 buffer[1183] = 18'b100000000000000000;
 buffer[1184] = 18'b100000000000000000;
 buffer[1185] = 18'b100000000000000000;
 buffer[1186] = 18'b100000000000000000;
 buffer[1187] = 18'b100000000000000000;
 buffer[1188] = 18'b100000000000000000;
 buffer[1189] = 18'b100000000000000000;
 buffer[1190] = 18'b100000000000000000;
 buffer[1191] = 18'b100000000000000000;
 buffer[1192] = 18'b100000000000000000;
 buffer[1193] = 18'b100000000000000000;
 buffer[1194] = 18'b100000000000000000;
 buffer[1195] = 18'b100000000000000000;
 buffer[1196] = 18'b100000000000000000;
 buffer[1197] = 18'b100000000000000000;
 buffer[1198] = 18'b100000000000000000;
 buffer[1199] = 18'b100000000000000000;
 buffer[1200] = 18'b100000000000000000;
 buffer[1201] = 18'b100000000000000000;
 buffer[1202] = 18'b100000000000000000;
 buffer[1203] = 18'b100000000000000000;
 buffer[1204] = 18'b100000000000000000;
 buffer[1205] = 18'b100000000000000000;
 buffer[1206] = 18'b100000000000000000;
 buffer[1207] = 18'b100000000000000000;
 buffer[1208] = 18'b100000000000000000;
 buffer[1209] = 18'b100000000000000000;
 buffer[1210] = 18'b100000000000000000;
 buffer[1211] = 18'b100000000000000000;
 buffer[1212] = 18'b100000000000000000;
 buffer[1213] = 18'b100000000000000000;
 buffer[1214] = 18'b100000000000000000;
 buffer[1215] = 18'b100000000000000000;
 buffer[1216] = 18'b100000000000000000;
 buffer[1217] = 18'b100000000000000000;
 buffer[1218] = 18'b100000000000000000;
 buffer[1219] = 18'b100000000000000000;
 buffer[1220] = 18'b100000000000000000;
 buffer[1221] = 18'b100000000000000000;
 buffer[1222] = 18'b100000000000000000;
 buffer[1223] = 18'b100000000000000000;
 buffer[1224] = 18'b100000000000000000;
 buffer[1225] = 18'b100000000000000000;
 buffer[1226] = 18'b100000000000000000;
 buffer[1227] = 18'b100000000000000000;
 buffer[1228] = 18'b100000000000000000;
 buffer[1229] = 18'b100000000000000000;
 buffer[1230] = 18'b100000000000000000;
 buffer[1231] = 18'b100000000000000000;
 buffer[1232] = 18'b100000000000000000;
 buffer[1233] = 18'b100000000000000000;
 buffer[1234] = 18'b100000000000000000;
 buffer[1235] = 18'b100000000000000000;
 buffer[1236] = 18'b100000000000000000;
 buffer[1237] = 18'b100000000000000000;
 buffer[1238] = 18'b100000000000000000;
 buffer[1239] = 18'b100000000000000000;
 buffer[1240] = 18'b100000000000000000;
 buffer[1241] = 18'b100000000000000000;
 buffer[1242] = 18'b100000000000000000;
 buffer[1243] = 18'b100000000000000000;
 buffer[1244] = 18'b100000000000000000;
 buffer[1245] = 18'b100000000000000000;
 buffer[1246] = 18'b100000000000000000;
 buffer[1247] = 18'b100000000000000000;
 buffer[1248] = 18'b100000000000000000;
 buffer[1249] = 18'b100000000000000000;
 buffer[1250] = 18'b100000000000000000;
 buffer[1251] = 18'b100000000000000000;
 buffer[1252] = 18'b100000000000000000;
 buffer[1253] = 18'b100000000000000000;
 buffer[1254] = 18'b100000000000000000;
 buffer[1255] = 18'b100000000000000000;
 buffer[1256] = 18'b100000000000000000;
 buffer[1257] = 18'b100000000000000000;
 buffer[1258] = 18'b100000000000000000;
 buffer[1259] = 18'b100000000000000000;
 buffer[1260] = 18'b100000000000000000;
 buffer[1261] = 18'b100000000000000000;
 buffer[1262] = 18'b100000000000000000;
 buffer[1263] = 18'b100000000000000000;
 buffer[1264] = 18'b100000000000000000;
 buffer[1265] = 18'b100000000000000000;
 buffer[1266] = 18'b100000000000000000;
 buffer[1267] = 18'b100000000000000000;
 buffer[1268] = 18'b100000000000000000;
 buffer[1269] = 18'b100000000000000000;
 buffer[1270] = 18'b100000000000000000;
 buffer[1271] = 18'b100000000000000000;
 buffer[1272] = 18'b100000000000000000;
 buffer[1273] = 18'b100000000000000000;
 buffer[1274] = 18'b100000000000000000;
 buffer[1275] = 18'b100000000000000000;
 buffer[1276] = 18'b100000000000000000;
 buffer[1277] = 18'b100000000000000000;
 buffer[1278] = 18'b100000000000000000;
 buffer[1279] = 18'b100000000000000000;
 buffer[1280] = 18'b100000000000000000;
 buffer[1281] = 18'b100000000000000000;
 buffer[1282] = 18'b100000000000000000;
 buffer[1283] = 18'b100000000000000000;
 buffer[1284] = 18'b100000000000000000;
 buffer[1285] = 18'b100000000000000000;
 buffer[1286] = 18'b100000000000000000;
 buffer[1287] = 18'b100000000000000000;
 buffer[1288] = 18'b100000000000000000;
 buffer[1289] = 18'b100000000000000000;
 buffer[1290] = 18'b100000000000000000;
 buffer[1291] = 18'b100000000000000000;
 buffer[1292] = 18'b100000000000000000;
 buffer[1293] = 18'b100000000000000000;
 buffer[1294] = 18'b100000000000000000;
 buffer[1295] = 18'b100000000000000000;
 buffer[1296] = 18'b100000000000000000;
 buffer[1297] = 18'b100000000000000000;
 buffer[1298] = 18'b100000000000000000;
 buffer[1299] = 18'b100000000000000000;
 buffer[1300] = 18'b100000000000000000;
 buffer[1301] = 18'b100000000000000000;
 buffer[1302] = 18'b100000000000000000;
 buffer[1303] = 18'b100000000000000000;
 buffer[1304] = 18'b100000000000000000;
 buffer[1305] = 18'b100000000000000000;
 buffer[1306] = 18'b100000000000000000;
 buffer[1307] = 18'b100000000000000000;
 buffer[1308] = 18'b100000000000000000;
 buffer[1309] = 18'b100000000000000000;
 buffer[1310] = 18'b100000000000000000;
 buffer[1311] = 18'b100000000000000000;
 buffer[1312] = 18'b100000000000000000;
 buffer[1313] = 18'b100000000000000000;
 buffer[1314] = 18'b100000000000000000;
 buffer[1315] = 18'b100000000000000000;
 buffer[1316] = 18'b100000000000000000;
 buffer[1317] = 18'b100000000000000000;
 buffer[1318] = 18'b100000000000000000;
 buffer[1319] = 18'b100000000000000000;
 buffer[1320] = 18'b100000000000000000;
 buffer[1321] = 18'b100000000000000000;
 buffer[1322] = 18'b100000000000000000;
 buffer[1323] = 18'b100000000000000000;
 buffer[1324] = 18'b100000000000000000;
 buffer[1325] = 18'b100000000000000000;
 buffer[1326] = 18'b100000000000000000;
 buffer[1327] = 18'b100000000000000000;
 buffer[1328] = 18'b100000000000000000;
 buffer[1329] = 18'b100000000000000000;
 buffer[1330] = 18'b100000000000000000;
 buffer[1331] = 18'b100000000000000000;
 buffer[1332] = 18'b100000000000000000;
 buffer[1333] = 18'b100000000000000000;
 buffer[1334] = 18'b100000000000000000;
 buffer[1335] = 18'b100000000000000000;
 buffer[1336] = 18'b100000000000000000;
 buffer[1337] = 18'b100000000000000000;
 buffer[1338] = 18'b100000000000000000;
 buffer[1339] = 18'b100000000000000000;
 buffer[1340] = 18'b100000000000000000;
 buffer[1341] = 18'b100000000000000000;
 buffer[1342] = 18'b100000000000000000;
 buffer[1343] = 18'b100000000000000000;
end

endmodule

module M_tilemap_mem_tiles_copy(
input      [10:0]                in_tiles_copy_addr0,
output reg  [17:0]     out_tiles_copy_rdata0,
output reg  [17:0]     out_tiles_copy_rdata1,
input      [0:0]             in_tiles_copy_wenable1,
input      [17:0]                 in_tiles_copy_wdata1,
input      [10:0]                in_tiles_copy_addr1,
input      clock0,
input      clock1
);
reg  [17:0] buffer[1343:0];
always @(posedge clock0) begin
  out_tiles_copy_rdata0 <= buffer[in_tiles_copy_addr0];
end
always @(posedge clock1) begin
  if (in_tiles_copy_wenable1) begin
    buffer[in_tiles_copy_addr1] <= in_tiles_copy_wdata1;
  end
end
initial begin
 buffer[0] = 18'b100000000000000000;
 buffer[1] = 18'b100000000000000000;
 buffer[2] = 18'b100000000000000000;
 buffer[3] = 18'b100000000000000000;
 buffer[4] = 18'b100000000000000000;
 buffer[5] = 18'b100000000000000000;
 buffer[6] = 18'b100000000000000000;
 buffer[7] = 18'b100000000000000000;
 buffer[8] = 18'b100000000000000000;
 buffer[9] = 18'b100000000000000000;
 buffer[10] = 18'b100000000000000000;
 buffer[11] = 18'b100000000000000000;
 buffer[12] = 18'b100000000000000000;
 buffer[13] = 18'b100000000000000000;
 buffer[14] = 18'b100000000000000000;
 buffer[15] = 18'b100000000000000000;
 buffer[16] = 18'b100000000000000000;
 buffer[17] = 18'b100000000000000000;
 buffer[18] = 18'b100000000000000000;
 buffer[19] = 18'b100000000000000000;
 buffer[20] = 18'b100000000000000000;
 buffer[21] = 18'b100000000000000000;
 buffer[22] = 18'b100000000000000000;
 buffer[23] = 18'b100000000000000000;
 buffer[24] = 18'b100000000000000000;
 buffer[25] = 18'b100000000000000000;
 buffer[26] = 18'b100000000000000000;
 buffer[27] = 18'b100000000000000000;
 buffer[28] = 18'b100000000000000000;
 buffer[29] = 18'b100000000000000000;
 buffer[30] = 18'b100000000000000000;
 buffer[31] = 18'b100000000000000000;
 buffer[32] = 18'b100000000000000000;
 buffer[33] = 18'b100000000000000000;
 buffer[34] = 18'b100000000000000000;
 buffer[35] = 18'b100000000000000000;
 buffer[36] = 18'b100000000000000000;
 buffer[37] = 18'b100000000000000000;
 buffer[38] = 18'b100000000000000000;
 buffer[39] = 18'b100000000000000000;
 buffer[40] = 18'b100000000000000000;
 buffer[41] = 18'b100000000000000000;
 buffer[42] = 18'b100000000000000000;
 buffer[43] = 18'b100000000000000000;
 buffer[44] = 18'b100000000000000000;
 buffer[45] = 18'b100000000000000000;
 buffer[46] = 18'b100000000000000000;
 buffer[47] = 18'b100000000000000000;
 buffer[48] = 18'b100000000000000000;
 buffer[49] = 18'b100000000000000000;
 buffer[50] = 18'b100000000000000000;
 buffer[51] = 18'b100000000000000000;
 buffer[52] = 18'b100000000000000000;
 buffer[53] = 18'b100000000000000000;
 buffer[54] = 18'b100000000000000000;
 buffer[55] = 18'b100000000000000000;
 buffer[56] = 18'b100000000000000000;
 buffer[57] = 18'b100000000000000000;
 buffer[58] = 18'b100000000000000000;
 buffer[59] = 18'b100000000000000000;
 buffer[60] = 18'b100000000000000000;
 buffer[61] = 18'b100000000000000000;
 buffer[62] = 18'b100000000000000000;
 buffer[63] = 18'b100000000000000000;
 buffer[64] = 18'b100000000000000000;
 buffer[65] = 18'b100000000000000000;
 buffer[66] = 18'b100000000000000000;
 buffer[67] = 18'b100000000000000000;
 buffer[68] = 18'b100000000000000000;
 buffer[69] = 18'b100000000000000000;
 buffer[70] = 18'b100000000000000000;
 buffer[71] = 18'b100000000000000000;
 buffer[72] = 18'b100000000000000000;
 buffer[73] = 18'b100000000000000000;
 buffer[74] = 18'b100000000000000000;
 buffer[75] = 18'b100000000000000000;
 buffer[76] = 18'b100000000000000000;
 buffer[77] = 18'b100000000000000000;
 buffer[78] = 18'b100000000000000000;
 buffer[79] = 18'b100000000000000000;
 buffer[80] = 18'b100000000000000000;
 buffer[81] = 18'b100000000000000000;
 buffer[82] = 18'b100000000000000000;
 buffer[83] = 18'b100000000000000000;
 buffer[84] = 18'b100000000000000000;
 buffer[85] = 18'b100000000000000000;
 buffer[86] = 18'b100000000000000000;
 buffer[87] = 18'b100000000000000000;
 buffer[88] = 18'b100000000000000000;
 buffer[89] = 18'b100000000000000000;
 buffer[90] = 18'b100000000000000000;
 buffer[91] = 18'b100000000000000000;
 buffer[92] = 18'b100000000000000000;
 buffer[93] = 18'b100000000000000000;
 buffer[94] = 18'b100000000000000000;
 buffer[95] = 18'b100000000000000000;
 buffer[96] = 18'b100000000000000000;
 buffer[97] = 18'b100000000000000000;
 buffer[98] = 18'b100000000000000000;
 buffer[99] = 18'b100000000000000000;
 buffer[100] = 18'b100000000000000000;
 buffer[101] = 18'b100000000000000000;
 buffer[102] = 18'b100000000000000000;
 buffer[103] = 18'b100000000000000000;
 buffer[104] = 18'b100000000000000000;
 buffer[105] = 18'b100000000000000000;
 buffer[106] = 18'b100000000000000000;
 buffer[107] = 18'b100000000000000000;
 buffer[108] = 18'b100000000000000000;
 buffer[109] = 18'b100000000000000000;
 buffer[110] = 18'b100000000000000000;
 buffer[111] = 18'b100000000000000000;
 buffer[112] = 18'b100000000000000000;
 buffer[113] = 18'b100000000000000000;
 buffer[114] = 18'b100000000000000000;
 buffer[115] = 18'b100000000000000000;
 buffer[116] = 18'b100000000000000000;
 buffer[117] = 18'b100000000000000000;
 buffer[118] = 18'b100000000000000000;
 buffer[119] = 18'b100000000000000000;
 buffer[120] = 18'b100000000000000000;
 buffer[121] = 18'b100000000000000000;
 buffer[122] = 18'b100000000000000000;
 buffer[123] = 18'b100000000000000000;
 buffer[124] = 18'b100000000000000000;
 buffer[125] = 18'b100000000000000000;
 buffer[126] = 18'b100000000000000000;
 buffer[127] = 18'b100000000000000000;
 buffer[128] = 18'b100000000000000000;
 buffer[129] = 18'b100000000000000000;
 buffer[130] = 18'b100000000000000000;
 buffer[131] = 18'b100000000000000000;
 buffer[132] = 18'b100000000000000000;
 buffer[133] = 18'b100000000000000000;
 buffer[134] = 18'b100000000000000000;
 buffer[135] = 18'b100000000000000000;
 buffer[136] = 18'b100000000000000000;
 buffer[137] = 18'b100000000000000000;
 buffer[138] = 18'b100000000000000000;
 buffer[139] = 18'b100000000000000000;
 buffer[140] = 18'b100000000000000000;
 buffer[141] = 18'b100000000000000000;
 buffer[142] = 18'b100000000000000000;
 buffer[143] = 18'b100000000000000000;
 buffer[144] = 18'b100000000000000000;
 buffer[145] = 18'b100000000000000000;
 buffer[146] = 18'b100000000000000000;
 buffer[147] = 18'b100000000000000000;
 buffer[148] = 18'b100000000000000000;
 buffer[149] = 18'b100000000000000000;
 buffer[150] = 18'b100000000000000000;
 buffer[151] = 18'b100000000000000000;
 buffer[152] = 18'b100000000000000000;
 buffer[153] = 18'b100000000000000000;
 buffer[154] = 18'b100000000000000000;
 buffer[155] = 18'b100000000000000000;
 buffer[156] = 18'b100000000000000000;
 buffer[157] = 18'b100000000000000000;
 buffer[158] = 18'b100000000000000000;
 buffer[159] = 18'b100000000000000000;
 buffer[160] = 18'b100000000000000000;
 buffer[161] = 18'b100000000000000000;
 buffer[162] = 18'b100000000000000000;
 buffer[163] = 18'b100000000000000000;
 buffer[164] = 18'b100000000000000000;
 buffer[165] = 18'b100000000000000000;
 buffer[166] = 18'b100000000000000000;
 buffer[167] = 18'b100000000000000000;
 buffer[168] = 18'b100000000000000000;
 buffer[169] = 18'b100000000000000000;
 buffer[170] = 18'b100000000000000000;
 buffer[171] = 18'b100000000000000000;
 buffer[172] = 18'b100000000000000000;
 buffer[173] = 18'b100000000000000000;
 buffer[174] = 18'b100000000000000000;
 buffer[175] = 18'b100000000000000000;
 buffer[176] = 18'b100000000000000000;
 buffer[177] = 18'b100000000000000000;
 buffer[178] = 18'b100000000000000000;
 buffer[179] = 18'b100000000000000000;
 buffer[180] = 18'b100000000000000000;
 buffer[181] = 18'b100000000000000000;
 buffer[182] = 18'b100000000000000000;
 buffer[183] = 18'b100000000000000000;
 buffer[184] = 18'b100000000000000000;
 buffer[185] = 18'b100000000000000000;
 buffer[186] = 18'b100000000000000000;
 buffer[187] = 18'b100000000000000000;
 buffer[188] = 18'b100000000000000000;
 buffer[189] = 18'b100000000000000000;
 buffer[190] = 18'b100000000000000000;
 buffer[191] = 18'b100000000000000000;
 buffer[192] = 18'b100000000000000000;
 buffer[193] = 18'b100000000000000000;
 buffer[194] = 18'b100000000000000000;
 buffer[195] = 18'b100000000000000000;
 buffer[196] = 18'b100000000000000000;
 buffer[197] = 18'b100000000000000000;
 buffer[198] = 18'b100000000000000000;
 buffer[199] = 18'b100000000000000000;
 buffer[200] = 18'b100000000000000000;
 buffer[201] = 18'b100000000000000000;
 buffer[202] = 18'b100000000000000000;
 buffer[203] = 18'b100000000000000000;
 buffer[204] = 18'b100000000000000000;
 buffer[205] = 18'b100000000000000000;
 buffer[206] = 18'b100000000000000000;
 buffer[207] = 18'b100000000000000000;
 buffer[208] = 18'b100000000000000000;
 buffer[209] = 18'b100000000000000000;
 buffer[210] = 18'b100000000000000000;
 buffer[211] = 18'b100000000000000000;
 buffer[212] = 18'b100000000000000000;
 buffer[213] = 18'b100000000000000000;
 buffer[214] = 18'b100000000000000000;
 buffer[215] = 18'b100000000000000000;
 buffer[216] = 18'b100000000000000000;
 buffer[217] = 18'b100000000000000000;
 buffer[218] = 18'b100000000000000000;
 buffer[219] = 18'b100000000000000000;
 buffer[220] = 18'b100000000000000000;
 buffer[221] = 18'b100000000000000000;
 buffer[222] = 18'b100000000000000000;
 buffer[223] = 18'b100000000000000000;
 buffer[224] = 18'b100000000000000000;
 buffer[225] = 18'b100000000000000000;
 buffer[226] = 18'b100000000000000000;
 buffer[227] = 18'b100000000000000000;
 buffer[228] = 18'b100000000000000000;
 buffer[229] = 18'b100000000000000000;
 buffer[230] = 18'b100000000000000000;
 buffer[231] = 18'b100000000000000000;
 buffer[232] = 18'b100000000000000000;
 buffer[233] = 18'b100000000000000000;
 buffer[234] = 18'b100000000000000000;
 buffer[235] = 18'b100000000000000000;
 buffer[236] = 18'b100000000000000000;
 buffer[237] = 18'b100000000000000000;
 buffer[238] = 18'b100000000000000000;
 buffer[239] = 18'b100000000000000000;
 buffer[240] = 18'b100000000000000000;
 buffer[241] = 18'b100000000000000000;
 buffer[242] = 18'b100000000000000000;
 buffer[243] = 18'b100000000000000000;
 buffer[244] = 18'b100000000000000000;
 buffer[245] = 18'b100000000000000000;
 buffer[246] = 18'b100000000000000000;
 buffer[247] = 18'b100000000000000000;
 buffer[248] = 18'b100000000000000000;
 buffer[249] = 18'b100000000000000000;
 buffer[250] = 18'b100000000000000000;
 buffer[251] = 18'b100000000000000000;
 buffer[252] = 18'b100000000000000000;
 buffer[253] = 18'b100000000000000000;
 buffer[254] = 18'b100000000000000000;
 buffer[255] = 18'b100000000000000000;
 buffer[256] = 18'b100000000000000000;
 buffer[257] = 18'b100000000000000000;
 buffer[258] = 18'b100000000000000000;
 buffer[259] = 18'b100000000000000000;
 buffer[260] = 18'b100000000000000000;
 buffer[261] = 18'b100000000000000000;
 buffer[262] = 18'b100000000000000000;
 buffer[263] = 18'b100000000000000000;
 buffer[264] = 18'b100000000000000000;
 buffer[265] = 18'b100000000000000000;
 buffer[266] = 18'b100000000000000000;
 buffer[267] = 18'b100000000000000000;
 buffer[268] = 18'b100000000000000000;
 buffer[269] = 18'b100000000000000000;
 buffer[270] = 18'b100000000000000000;
 buffer[271] = 18'b100000000000000000;
 buffer[272] = 18'b100000000000000000;
 buffer[273] = 18'b100000000000000000;
 buffer[274] = 18'b100000000000000000;
 buffer[275] = 18'b100000000000000000;
 buffer[276] = 18'b100000000000000000;
 buffer[277] = 18'b100000000000000000;
 buffer[278] = 18'b100000000000000000;
 buffer[279] = 18'b100000000000000000;
 buffer[280] = 18'b100000000000000000;
 buffer[281] = 18'b100000000000000000;
 buffer[282] = 18'b100000000000000000;
 buffer[283] = 18'b100000000000000000;
 buffer[284] = 18'b100000000000000000;
 buffer[285] = 18'b100000000000000000;
 buffer[286] = 18'b100000000000000000;
 buffer[287] = 18'b100000000000000000;
 buffer[288] = 18'b100000000000000000;
 buffer[289] = 18'b100000000000000000;
 buffer[290] = 18'b100000000000000000;
 buffer[291] = 18'b100000000000000000;
 buffer[292] = 18'b100000000000000000;
 buffer[293] = 18'b100000000000000000;
 buffer[294] = 18'b100000000000000000;
 buffer[295] = 18'b100000000000000000;
 buffer[296] = 18'b100000000000000000;
 buffer[297] = 18'b100000000000000000;
 buffer[298] = 18'b100000000000000000;
 buffer[299] = 18'b100000000000000000;
 buffer[300] = 18'b100000000000000000;
 buffer[301] = 18'b100000000000000000;
 buffer[302] = 18'b100000000000000000;
 buffer[303] = 18'b100000000000000000;
 buffer[304] = 18'b100000000000000000;
 buffer[305] = 18'b100000000000000000;
 buffer[306] = 18'b100000000000000000;
 buffer[307] = 18'b100000000000000000;
 buffer[308] = 18'b100000000000000000;
 buffer[309] = 18'b100000000000000000;
 buffer[310] = 18'b100000000000000000;
 buffer[311] = 18'b100000000000000000;
 buffer[312] = 18'b100000000000000000;
 buffer[313] = 18'b100000000000000000;
 buffer[314] = 18'b100000000000000000;
 buffer[315] = 18'b100000000000000000;
 buffer[316] = 18'b100000000000000000;
 buffer[317] = 18'b100000000000000000;
 buffer[318] = 18'b100000000000000000;
 buffer[319] = 18'b100000000000000000;
 buffer[320] = 18'b100000000000000000;
 buffer[321] = 18'b100000000000000000;
 buffer[322] = 18'b100000000000000000;
 buffer[323] = 18'b100000000000000000;
 buffer[324] = 18'b100000000000000000;
 buffer[325] = 18'b100000000000000000;
 buffer[326] = 18'b100000000000000000;
 buffer[327] = 18'b100000000000000000;
 buffer[328] = 18'b100000000000000000;
 buffer[329] = 18'b100000000000000000;
 buffer[330] = 18'b100000000000000000;
 buffer[331] = 18'b100000000000000000;
 buffer[332] = 18'b100000000000000000;
 buffer[333] = 18'b100000000000000000;
 buffer[334] = 18'b100000000000000000;
 buffer[335] = 18'b100000000000000000;
 buffer[336] = 18'b100000000000000000;
 buffer[337] = 18'b100000000000000000;
 buffer[338] = 18'b100000000000000000;
 buffer[339] = 18'b100000000000000000;
 buffer[340] = 18'b100000000000000000;
 buffer[341] = 18'b100000000000000000;
 buffer[342] = 18'b100000000000000000;
 buffer[343] = 18'b100000000000000000;
 buffer[344] = 18'b100000000000000000;
 buffer[345] = 18'b100000000000000000;
 buffer[346] = 18'b100000000000000000;
 buffer[347] = 18'b100000000000000000;
 buffer[348] = 18'b100000000000000000;
 buffer[349] = 18'b100000000000000000;
 buffer[350] = 18'b100000000000000000;
 buffer[351] = 18'b100000000000000000;
 buffer[352] = 18'b100000000000000000;
 buffer[353] = 18'b100000000000000000;
 buffer[354] = 18'b100000000000000000;
 buffer[355] = 18'b100000000000000000;
 buffer[356] = 18'b100000000000000000;
 buffer[357] = 18'b100000000000000000;
 buffer[358] = 18'b100000000000000000;
 buffer[359] = 18'b100000000000000000;
 buffer[360] = 18'b100000000000000000;
 buffer[361] = 18'b100000000000000000;
 buffer[362] = 18'b100000000000000000;
 buffer[363] = 18'b100000000000000000;
 buffer[364] = 18'b100000000000000000;
 buffer[365] = 18'b100000000000000000;
 buffer[366] = 18'b100000000000000000;
 buffer[367] = 18'b100000000000000000;
 buffer[368] = 18'b100000000000000000;
 buffer[369] = 18'b100000000000000000;
 buffer[370] = 18'b100000000000000000;
 buffer[371] = 18'b100000000000000000;
 buffer[372] = 18'b100000000000000000;
 buffer[373] = 18'b100000000000000000;
 buffer[374] = 18'b100000000000000000;
 buffer[375] = 18'b100000000000000000;
 buffer[376] = 18'b100000000000000000;
 buffer[377] = 18'b100000000000000000;
 buffer[378] = 18'b100000000000000000;
 buffer[379] = 18'b100000000000000000;
 buffer[380] = 18'b100000000000000000;
 buffer[381] = 18'b100000000000000000;
 buffer[382] = 18'b100000000000000000;
 buffer[383] = 18'b100000000000000000;
 buffer[384] = 18'b100000000000000000;
 buffer[385] = 18'b100000000000000000;
 buffer[386] = 18'b100000000000000000;
 buffer[387] = 18'b100000000000000000;
 buffer[388] = 18'b100000000000000000;
 buffer[389] = 18'b100000000000000000;
 buffer[390] = 18'b100000000000000000;
 buffer[391] = 18'b100000000000000000;
 buffer[392] = 18'b100000000000000000;
 buffer[393] = 18'b100000000000000000;
 buffer[394] = 18'b100000000000000000;
 buffer[395] = 18'b100000000000000000;
 buffer[396] = 18'b100000000000000000;
 buffer[397] = 18'b100000000000000000;
 buffer[398] = 18'b100000000000000000;
 buffer[399] = 18'b100000000000000000;
 buffer[400] = 18'b100000000000000000;
 buffer[401] = 18'b100000000000000000;
 buffer[402] = 18'b100000000000000000;
 buffer[403] = 18'b100000000000000000;
 buffer[404] = 18'b100000000000000000;
 buffer[405] = 18'b100000000000000000;
 buffer[406] = 18'b100000000000000000;
 buffer[407] = 18'b100000000000000000;
 buffer[408] = 18'b100000000000000000;
 buffer[409] = 18'b100000000000000000;
 buffer[410] = 18'b100000000000000000;
 buffer[411] = 18'b100000000000000000;
 buffer[412] = 18'b100000000000000000;
 buffer[413] = 18'b100000000000000000;
 buffer[414] = 18'b100000000000000000;
 buffer[415] = 18'b100000000000000000;
 buffer[416] = 18'b100000000000000000;
 buffer[417] = 18'b100000000000000000;
 buffer[418] = 18'b100000000000000000;
 buffer[419] = 18'b100000000000000000;
 buffer[420] = 18'b100000000000000000;
 buffer[421] = 18'b100000000000000000;
 buffer[422] = 18'b100000000000000000;
 buffer[423] = 18'b100000000000000000;
 buffer[424] = 18'b100000000000000000;
 buffer[425] = 18'b100000000000000000;
 buffer[426] = 18'b100000000000000000;
 buffer[427] = 18'b100000000000000000;
 buffer[428] = 18'b100000000000000000;
 buffer[429] = 18'b100000000000000000;
 buffer[430] = 18'b100000000000000000;
 buffer[431] = 18'b100000000000000000;
 buffer[432] = 18'b100000000000000000;
 buffer[433] = 18'b100000000000000000;
 buffer[434] = 18'b100000000000000000;
 buffer[435] = 18'b100000000000000000;
 buffer[436] = 18'b100000000000000000;
 buffer[437] = 18'b100000000000000000;
 buffer[438] = 18'b100000000000000000;
 buffer[439] = 18'b100000000000000000;
 buffer[440] = 18'b100000000000000000;
 buffer[441] = 18'b100000000000000000;
 buffer[442] = 18'b100000000000000000;
 buffer[443] = 18'b100000000000000000;
 buffer[444] = 18'b100000000000000000;
 buffer[445] = 18'b100000000000000000;
 buffer[446] = 18'b100000000000000000;
 buffer[447] = 18'b100000000000000000;
 buffer[448] = 18'b100000000000000000;
 buffer[449] = 18'b100000000000000000;
 buffer[450] = 18'b100000000000000000;
 buffer[451] = 18'b100000000000000000;
 buffer[452] = 18'b100000000000000000;
 buffer[453] = 18'b100000000000000000;
 buffer[454] = 18'b100000000000000000;
 buffer[455] = 18'b100000000000000000;
 buffer[456] = 18'b100000000000000000;
 buffer[457] = 18'b100000000000000000;
 buffer[458] = 18'b100000000000000000;
 buffer[459] = 18'b100000000000000000;
 buffer[460] = 18'b100000000000000000;
 buffer[461] = 18'b100000000000000000;
 buffer[462] = 18'b100000000000000000;
 buffer[463] = 18'b100000000000000000;
 buffer[464] = 18'b100000000000000000;
 buffer[465] = 18'b100000000000000000;
 buffer[466] = 18'b100000000000000000;
 buffer[467] = 18'b100000000000000000;
 buffer[468] = 18'b100000000000000000;
 buffer[469] = 18'b100000000000000000;
 buffer[470] = 18'b100000000000000000;
 buffer[471] = 18'b100000000000000000;
 buffer[472] = 18'b100000000000000000;
 buffer[473] = 18'b100000000000000000;
 buffer[474] = 18'b100000000000000000;
 buffer[475] = 18'b100000000000000000;
 buffer[476] = 18'b100000000000000000;
 buffer[477] = 18'b100000000000000000;
 buffer[478] = 18'b100000000000000000;
 buffer[479] = 18'b100000000000000000;
 buffer[480] = 18'b100000000000000000;
 buffer[481] = 18'b100000000000000000;
 buffer[482] = 18'b100000000000000000;
 buffer[483] = 18'b100000000000000000;
 buffer[484] = 18'b100000000000000000;
 buffer[485] = 18'b100000000000000000;
 buffer[486] = 18'b100000000000000000;
 buffer[487] = 18'b100000000000000000;
 buffer[488] = 18'b100000000000000000;
 buffer[489] = 18'b100000000000000000;
 buffer[490] = 18'b100000000000000000;
 buffer[491] = 18'b100000000000000000;
 buffer[492] = 18'b100000000000000000;
 buffer[493] = 18'b100000000000000000;
 buffer[494] = 18'b100000000000000000;
 buffer[495] = 18'b100000000000000000;
 buffer[496] = 18'b100000000000000000;
 buffer[497] = 18'b100000000000000000;
 buffer[498] = 18'b100000000000000000;
 buffer[499] = 18'b100000000000000000;
 buffer[500] = 18'b100000000000000000;
 buffer[501] = 18'b100000000000000000;
 buffer[502] = 18'b100000000000000000;
 buffer[503] = 18'b100000000000000000;
 buffer[504] = 18'b100000000000000000;
 buffer[505] = 18'b100000000000000000;
 buffer[506] = 18'b100000000000000000;
 buffer[507] = 18'b100000000000000000;
 buffer[508] = 18'b100000000000000000;
 buffer[509] = 18'b100000000000000000;
 buffer[510] = 18'b100000000000000000;
 buffer[511] = 18'b100000000000000000;
 buffer[512] = 18'b100000000000000000;
 buffer[513] = 18'b100000000000000000;
 buffer[514] = 18'b100000000000000000;
 buffer[515] = 18'b100000000000000000;
 buffer[516] = 18'b100000000000000000;
 buffer[517] = 18'b100000000000000000;
 buffer[518] = 18'b100000000000000000;
 buffer[519] = 18'b100000000000000000;
 buffer[520] = 18'b100000000000000000;
 buffer[521] = 18'b100000000000000000;
 buffer[522] = 18'b100000000000000000;
 buffer[523] = 18'b100000000000000000;
 buffer[524] = 18'b100000000000000000;
 buffer[525] = 18'b100000000000000000;
 buffer[526] = 18'b100000000000000000;
 buffer[527] = 18'b100000000000000000;
 buffer[528] = 18'b100000000000000000;
 buffer[529] = 18'b100000000000000000;
 buffer[530] = 18'b100000000000000000;
 buffer[531] = 18'b100000000000000000;
 buffer[532] = 18'b100000000000000000;
 buffer[533] = 18'b100000000000000000;
 buffer[534] = 18'b100000000000000000;
 buffer[535] = 18'b100000000000000000;
 buffer[536] = 18'b100000000000000000;
 buffer[537] = 18'b100000000000000000;
 buffer[538] = 18'b100000000000000000;
 buffer[539] = 18'b100000000000000000;
 buffer[540] = 18'b100000000000000000;
 buffer[541] = 18'b100000000000000000;
 buffer[542] = 18'b100000000000000000;
 buffer[543] = 18'b100000000000000000;
 buffer[544] = 18'b100000000000000000;
 buffer[545] = 18'b100000000000000000;
 buffer[546] = 18'b100000000000000000;
 buffer[547] = 18'b100000000000000000;
 buffer[548] = 18'b100000000000000000;
 buffer[549] = 18'b100000000000000000;
 buffer[550] = 18'b100000000000000000;
 buffer[551] = 18'b100000000000000000;
 buffer[552] = 18'b100000000000000000;
 buffer[553] = 18'b100000000000000000;
 buffer[554] = 18'b100000000000000000;
 buffer[555] = 18'b100000000000000000;
 buffer[556] = 18'b100000000000000000;
 buffer[557] = 18'b100000000000000000;
 buffer[558] = 18'b100000000000000000;
 buffer[559] = 18'b100000000000000000;
 buffer[560] = 18'b100000000000000000;
 buffer[561] = 18'b100000000000000000;
 buffer[562] = 18'b100000000000000000;
 buffer[563] = 18'b100000000000000000;
 buffer[564] = 18'b100000000000000000;
 buffer[565] = 18'b100000000000000000;
 buffer[566] = 18'b100000000000000000;
 buffer[567] = 18'b100000000000000000;
 buffer[568] = 18'b100000000000000000;
 buffer[569] = 18'b100000000000000000;
 buffer[570] = 18'b100000000000000000;
 buffer[571] = 18'b100000000000000000;
 buffer[572] = 18'b100000000000000000;
 buffer[573] = 18'b100000000000000000;
 buffer[574] = 18'b100000000000000000;
 buffer[575] = 18'b100000000000000000;
 buffer[576] = 18'b100000000000000000;
 buffer[577] = 18'b100000000000000000;
 buffer[578] = 18'b100000000000000000;
 buffer[579] = 18'b100000000000000000;
 buffer[580] = 18'b100000000000000000;
 buffer[581] = 18'b100000000000000000;
 buffer[582] = 18'b100000000000000000;
 buffer[583] = 18'b100000000000000000;
 buffer[584] = 18'b100000000000000000;
 buffer[585] = 18'b100000000000000000;
 buffer[586] = 18'b100000000000000000;
 buffer[587] = 18'b100000000000000000;
 buffer[588] = 18'b100000000000000000;
 buffer[589] = 18'b100000000000000000;
 buffer[590] = 18'b100000000000000000;
 buffer[591] = 18'b100000000000000000;
 buffer[592] = 18'b100000000000000000;
 buffer[593] = 18'b100000000000000000;
 buffer[594] = 18'b100000000000000000;
 buffer[595] = 18'b100000000000000000;
 buffer[596] = 18'b100000000000000000;
 buffer[597] = 18'b100000000000000000;
 buffer[598] = 18'b100000000000000000;
 buffer[599] = 18'b100000000000000000;
 buffer[600] = 18'b100000000000000000;
 buffer[601] = 18'b100000000000000000;
 buffer[602] = 18'b100000000000000000;
 buffer[603] = 18'b100000000000000000;
 buffer[604] = 18'b100000000000000000;
 buffer[605] = 18'b100000000000000000;
 buffer[606] = 18'b100000000000000000;
 buffer[607] = 18'b100000000000000000;
 buffer[608] = 18'b100000000000000000;
 buffer[609] = 18'b100000000000000000;
 buffer[610] = 18'b100000000000000000;
 buffer[611] = 18'b100000000000000000;
 buffer[612] = 18'b100000000000000000;
 buffer[613] = 18'b100000000000000000;
 buffer[614] = 18'b100000000000000000;
 buffer[615] = 18'b100000000000000000;
 buffer[616] = 18'b100000000000000000;
 buffer[617] = 18'b100000000000000000;
 buffer[618] = 18'b100000000000000000;
 buffer[619] = 18'b100000000000000000;
 buffer[620] = 18'b100000000000000000;
 buffer[621] = 18'b100000000000000000;
 buffer[622] = 18'b100000000000000000;
 buffer[623] = 18'b100000000000000000;
 buffer[624] = 18'b100000000000000000;
 buffer[625] = 18'b100000000000000000;
 buffer[626] = 18'b100000000000000000;
 buffer[627] = 18'b100000000000000000;
 buffer[628] = 18'b100000000000000000;
 buffer[629] = 18'b100000000000000000;
 buffer[630] = 18'b100000000000000000;
 buffer[631] = 18'b100000000000000000;
 buffer[632] = 18'b100000000000000000;
 buffer[633] = 18'b100000000000000000;
 buffer[634] = 18'b100000000000000000;
 buffer[635] = 18'b100000000000000000;
 buffer[636] = 18'b100000000000000000;
 buffer[637] = 18'b100000000000000000;
 buffer[638] = 18'b100000000000000000;
 buffer[639] = 18'b100000000000000000;
 buffer[640] = 18'b100000000000000000;
 buffer[641] = 18'b100000000000000000;
 buffer[642] = 18'b100000000000000000;
 buffer[643] = 18'b100000000000000000;
 buffer[644] = 18'b100000000000000000;
 buffer[645] = 18'b100000000000000000;
 buffer[646] = 18'b100000000000000000;
 buffer[647] = 18'b100000000000000000;
 buffer[648] = 18'b100000000000000000;
 buffer[649] = 18'b100000000000000000;
 buffer[650] = 18'b100000000000000000;
 buffer[651] = 18'b100000000000000000;
 buffer[652] = 18'b100000000000000000;
 buffer[653] = 18'b100000000000000000;
 buffer[654] = 18'b100000000000000000;
 buffer[655] = 18'b100000000000000000;
 buffer[656] = 18'b100000000000000000;
 buffer[657] = 18'b100000000000000000;
 buffer[658] = 18'b100000000000000000;
 buffer[659] = 18'b100000000000000000;
 buffer[660] = 18'b100000000000000000;
 buffer[661] = 18'b100000000000000000;
 buffer[662] = 18'b100000000000000000;
 buffer[663] = 18'b100000000000000000;
 buffer[664] = 18'b100000000000000000;
 buffer[665] = 18'b100000000000000000;
 buffer[666] = 18'b100000000000000000;
 buffer[667] = 18'b100000000000000000;
 buffer[668] = 18'b100000000000000000;
 buffer[669] = 18'b100000000000000000;
 buffer[670] = 18'b100000000000000000;
 buffer[671] = 18'b100000000000000000;
 buffer[672] = 18'b100000000000000000;
 buffer[673] = 18'b100000000000000000;
 buffer[674] = 18'b100000000000000000;
 buffer[675] = 18'b100000000000000000;
 buffer[676] = 18'b100000000000000000;
 buffer[677] = 18'b100000000000000000;
 buffer[678] = 18'b100000000000000000;
 buffer[679] = 18'b100000000000000000;
 buffer[680] = 18'b100000000000000000;
 buffer[681] = 18'b100000000000000000;
 buffer[682] = 18'b100000000000000000;
 buffer[683] = 18'b100000000000000000;
 buffer[684] = 18'b100000000000000000;
 buffer[685] = 18'b100000000000000000;
 buffer[686] = 18'b100000000000000000;
 buffer[687] = 18'b100000000000000000;
 buffer[688] = 18'b100000000000000000;
 buffer[689] = 18'b100000000000000000;
 buffer[690] = 18'b100000000000000000;
 buffer[691] = 18'b100000000000000000;
 buffer[692] = 18'b100000000000000000;
 buffer[693] = 18'b100000000000000000;
 buffer[694] = 18'b100000000000000000;
 buffer[695] = 18'b100000000000000000;
 buffer[696] = 18'b100000000000000000;
 buffer[697] = 18'b100000000000000000;
 buffer[698] = 18'b100000000000000000;
 buffer[699] = 18'b100000000000000000;
 buffer[700] = 18'b100000000000000000;
 buffer[701] = 18'b100000000000000000;
 buffer[702] = 18'b100000000000000000;
 buffer[703] = 18'b100000000000000000;
 buffer[704] = 18'b100000000000000000;
 buffer[705] = 18'b100000000000000000;
 buffer[706] = 18'b100000000000000000;
 buffer[707] = 18'b100000000000000000;
 buffer[708] = 18'b100000000000000000;
 buffer[709] = 18'b100000000000000000;
 buffer[710] = 18'b100000000000000000;
 buffer[711] = 18'b100000000000000000;
 buffer[712] = 18'b100000000000000000;
 buffer[713] = 18'b100000000000000000;
 buffer[714] = 18'b100000000000000000;
 buffer[715] = 18'b100000000000000000;
 buffer[716] = 18'b100000000000000000;
 buffer[717] = 18'b100000000000000000;
 buffer[718] = 18'b100000000000000000;
 buffer[719] = 18'b100000000000000000;
 buffer[720] = 18'b100000000000000000;
 buffer[721] = 18'b100000000000000000;
 buffer[722] = 18'b100000000000000000;
 buffer[723] = 18'b100000000000000000;
 buffer[724] = 18'b100000000000000000;
 buffer[725] = 18'b100000000000000000;
 buffer[726] = 18'b100000000000000000;
 buffer[727] = 18'b100000000000000000;
 buffer[728] = 18'b100000000000000000;
 buffer[729] = 18'b100000000000000000;
 buffer[730] = 18'b100000000000000000;
 buffer[731] = 18'b100000000000000000;
 buffer[732] = 18'b100000000000000000;
 buffer[733] = 18'b100000000000000000;
 buffer[734] = 18'b100000000000000000;
 buffer[735] = 18'b100000000000000000;
 buffer[736] = 18'b100000000000000000;
 buffer[737] = 18'b100000000000000000;
 buffer[738] = 18'b100000000000000000;
 buffer[739] = 18'b100000000000000000;
 buffer[740] = 18'b100000000000000000;
 buffer[741] = 18'b100000000000000000;
 buffer[742] = 18'b100000000000000000;
 buffer[743] = 18'b100000000000000000;
 buffer[744] = 18'b100000000000000000;
 buffer[745] = 18'b100000000000000000;
 buffer[746] = 18'b100000000000000000;
 buffer[747] = 18'b100000000000000000;
 buffer[748] = 18'b100000000000000000;
 buffer[749] = 18'b100000000000000000;
 buffer[750] = 18'b100000000000000000;
 buffer[751] = 18'b100000000000000000;
 buffer[752] = 18'b100000000000000000;
 buffer[753] = 18'b100000000000000000;
 buffer[754] = 18'b100000000000000000;
 buffer[755] = 18'b100000000000000000;
 buffer[756] = 18'b100000000000000000;
 buffer[757] = 18'b100000000000000000;
 buffer[758] = 18'b100000000000000000;
 buffer[759] = 18'b100000000000000000;
 buffer[760] = 18'b100000000000000000;
 buffer[761] = 18'b100000000000000000;
 buffer[762] = 18'b100000000000000000;
 buffer[763] = 18'b100000000000000000;
 buffer[764] = 18'b100000000000000000;
 buffer[765] = 18'b100000000000000000;
 buffer[766] = 18'b100000000000000000;
 buffer[767] = 18'b100000000000000000;
 buffer[768] = 18'b100000000000000000;
 buffer[769] = 18'b100000000000000000;
 buffer[770] = 18'b100000000000000000;
 buffer[771] = 18'b100000000000000000;
 buffer[772] = 18'b100000000000000000;
 buffer[773] = 18'b100000000000000000;
 buffer[774] = 18'b100000000000000000;
 buffer[775] = 18'b100000000000000000;
 buffer[776] = 18'b100000000000000000;
 buffer[777] = 18'b100000000000000000;
 buffer[778] = 18'b100000000000000000;
 buffer[779] = 18'b100000000000000000;
 buffer[780] = 18'b100000000000000000;
 buffer[781] = 18'b100000000000000000;
 buffer[782] = 18'b100000000000000000;
 buffer[783] = 18'b100000000000000000;
 buffer[784] = 18'b100000000000000000;
 buffer[785] = 18'b100000000000000000;
 buffer[786] = 18'b100000000000000000;
 buffer[787] = 18'b100000000000000000;
 buffer[788] = 18'b100000000000000000;
 buffer[789] = 18'b100000000000000000;
 buffer[790] = 18'b100000000000000000;
 buffer[791] = 18'b100000000000000000;
 buffer[792] = 18'b100000000000000000;
 buffer[793] = 18'b100000000000000000;
 buffer[794] = 18'b100000000000000000;
 buffer[795] = 18'b100000000000000000;
 buffer[796] = 18'b100000000000000000;
 buffer[797] = 18'b100000000000000000;
 buffer[798] = 18'b100000000000000000;
 buffer[799] = 18'b100000000000000000;
 buffer[800] = 18'b100000000000000000;
 buffer[801] = 18'b100000000000000000;
 buffer[802] = 18'b100000000000000000;
 buffer[803] = 18'b100000000000000000;
 buffer[804] = 18'b100000000000000000;
 buffer[805] = 18'b100000000000000000;
 buffer[806] = 18'b100000000000000000;
 buffer[807] = 18'b100000000000000000;
 buffer[808] = 18'b100000000000000000;
 buffer[809] = 18'b100000000000000000;
 buffer[810] = 18'b100000000000000000;
 buffer[811] = 18'b100000000000000000;
 buffer[812] = 18'b100000000000000000;
 buffer[813] = 18'b100000000000000000;
 buffer[814] = 18'b100000000000000000;
 buffer[815] = 18'b100000000000000000;
 buffer[816] = 18'b100000000000000000;
 buffer[817] = 18'b100000000000000000;
 buffer[818] = 18'b100000000000000000;
 buffer[819] = 18'b100000000000000000;
 buffer[820] = 18'b100000000000000000;
 buffer[821] = 18'b100000000000000000;
 buffer[822] = 18'b100000000000000000;
 buffer[823] = 18'b100000000000000000;
 buffer[824] = 18'b100000000000000000;
 buffer[825] = 18'b100000000000000000;
 buffer[826] = 18'b100000000000000000;
 buffer[827] = 18'b100000000000000000;
 buffer[828] = 18'b100000000000000000;
 buffer[829] = 18'b100000000000000000;
 buffer[830] = 18'b100000000000000000;
 buffer[831] = 18'b100000000000000000;
 buffer[832] = 18'b100000000000000000;
 buffer[833] = 18'b100000000000000000;
 buffer[834] = 18'b100000000000000000;
 buffer[835] = 18'b100000000000000000;
 buffer[836] = 18'b100000000000000000;
 buffer[837] = 18'b100000000000000000;
 buffer[838] = 18'b100000000000000000;
 buffer[839] = 18'b100000000000000000;
 buffer[840] = 18'b100000000000000000;
 buffer[841] = 18'b100000000000000000;
 buffer[842] = 18'b100000000000000000;
 buffer[843] = 18'b100000000000000000;
 buffer[844] = 18'b100000000000000000;
 buffer[845] = 18'b100000000000000000;
 buffer[846] = 18'b100000000000000000;
 buffer[847] = 18'b100000000000000000;
 buffer[848] = 18'b100000000000000000;
 buffer[849] = 18'b100000000000000000;
 buffer[850] = 18'b100000000000000000;
 buffer[851] = 18'b100000000000000000;
 buffer[852] = 18'b100000000000000000;
 buffer[853] = 18'b100000000000000000;
 buffer[854] = 18'b100000000000000000;
 buffer[855] = 18'b100000000000000000;
 buffer[856] = 18'b100000000000000000;
 buffer[857] = 18'b100000000000000000;
 buffer[858] = 18'b100000000000000000;
 buffer[859] = 18'b100000000000000000;
 buffer[860] = 18'b100000000000000000;
 buffer[861] = 18'b100000000000000000;
 buffer[862] = 18'b100000000000000000;
 buffer[863] = 18'b100000000000000000;
 buffer[864] = 18'b100000000000000000;
 buffer[865] = 18'b100000000000000000;
 buffer[866] = 18'b100000000000000000;
 buffer[867] = 18'b100000000000000000;
 buffer[868] = 18'b100000000000000000;
 buffer[869] = 18'b100000000000000000;
 buffer[870] = 18'b100000000000000000;
 buffer[871] = 18'b100000000000000000;
 buffer[872] = 18'b100000000000000000;
 buffer[873] = 18'b100000000000000000;
 buffer[874] = 18'b100000000000000000;
 buffer[875] = 18'b100000000000000000;
 buffer[876] = 18'b100000000000000000;
 buffer[877] = 18'b100000000000000000;
 buffer[878] = 18'b100000000000000000;
 buffer[879] = 18'b100000000000000000;
 buffer[880] = 18'b100000000000000000;
 buffer[881] = 18'b100000000000000000;
 buffer[882] = 18'b100000000000000000;
 buffer[883] = 18'b100000000000000000;
 buffer[884] = 18'b100000000000000000;
 buffer[885] = 18'b100000000000000000;
 buffer[886] = 18'b100000000000000000;
 buffer[887] = 18'b100000000000000000;
 buffer[888] = 18'b100000000000000000;
 buffer[889] = 18'b100000000000000000;
 buffer[890] = 18'b100000000000000000;
 buffer[891] = 18'b100000000000000000;
 buffer[892] = 18'b100000000000000000;
 buffer[893] = 18'b100000000000000000;
 buffer[894] = 18'b100000000000000000;
 buffer[895] = 18'b100000000000000000;
 buffer[896] = 18'b100000000000000000;
 buffer[897] = 18'b100000000000000000;
 buffer[898] = 18'b100000000000000000;
 buffer[899] = 18'b100000000000000000;
 buffer[900] = 18'b100000000000000000;
 buffer[901] = 18'b100000000000000000;
 buffer[902] = 18'b100000000000000000;
 buffer[903] = 18'b100000000000000000;
 buffer[904] = 18'b100000000000000000;
 buffer[905] = 18'b100000000000000000;
 buffer[906] = 18'b100000000000000000;
 buffer[907] = 18'b100000000000000000;
 buffer[908] = 18'b100000000000000000;
 buffer[909] = 18'b100000000000000000;
 buffer[910] = 18'b100000000000000000;
 buffer[911] = 18'b100000000000000000;
 buffer[912] = 18'b100000000000000000;
 buffer[913] = 18'b100000000000000000;
 buffer[914] = 18'b100000000000000000;
 buffer[915] = 18'b100000000000000000;
 buffer[916] = 18'b100000000000000000;
 buffer[917] = 18'b100000000000000000;
 buffer[918] = 18'b100000000000000000;
 buffer[919] = 18'b100000000000000000;
 buffer[920] = 18'b100000000000000000;
 buffer[921] = 18'b100000000000000000;
 buffer[922] = 18'b100000000000000000;
 buffer[923] = 18'b100000000000000000;
 buffer[924] = 18'b100000000000000000;
 buffer[925] = 18'b100000000000000000;
 buffer[926] = 18'b100000000000000000;
 buffer[927] = 18'b100000000000000000;
 buffer[928] = 18'b100000000000000000;
 buffer[929] = 18'b100000000000000000;
 buffer[930] = 18'b100000000000000000;
 buffer[931] = 18'b100000000000000000;
 buffer[932] = 18'b100000000000000000;
 buffer[933] = 18'b100000000000000000;
 buffer[934] = 18'b100000000000000000;
 buffer[935] = 18'b100000000000000000;
 buffer[936] = 18'b100000000000000000;
 buffer[937] = 18'b100000000000000000;
 buffer[938] = 18'b100000000000000000;
 buffer[939] = 18'b100000000000000000;
 buffer[940] = 18'b100000000000000000;
 buffer[941] = 18'b100000000000000000;
 buffer[942] = 18'b100000000000000000;
 buffer[943] = 18'b100000000000000000;
 buffer[944] = 18'b100000000000000000;
 buffer[945] = 18'b100000000000000000;
 buffer[946] = 18'b100000000000000000;
 buffer[947] = 18'b100000000000000000;
 buffer[948] = 18'b100000000000000000;
 buffer[949] = 18'b100000000000000000;
 buffer[950] = 18'b100000000000000000;
 buffer[951] = 18'b100000000000000000;
 buffer[952] = 18'b100000000000000000;
 buffer[953] = 18'b100000000000000000;
 buffer[954] = 18'b100000000000000000;
 buffer[955] = 18'b100000000000000000;
 buffer[956] = 18'b100000000000000000;
 buffer[957] = 18'b100000000000000000;
 buffer[958] = 18'b100000000000000000;
 buffer[959] = 18'b100000000000000000;
 buffer[960] = 18'b100000000000000000;
 buffer[961] = 18'b100000000000000000;
 buffer[962] = 18'b100000000000000000;
 buffer[963] = 18'b100000000000000000;
 buffer[964] = 18'b100000000000000000;
 buffer[965] = 18'b100000000000000000;
 buffer[966] = 18'b100000000000000000;
 buffer[967] = 18'b100000000000000000;
 buffer[968] = 18'b100000000000000000;
 buffer[969] = 18'b100000000000000000;
 buffer[970] = 18'b100000000000000000;
 buffer[971] = 18'b100000000000000000;
 buffer[972] = 18'b100000000000000000;
 buffer[973] = 18'b100000000000000000;
 buffer[974] = 18'b100000000000000000;
 buffer[975] = 18'b100000000000000000;
 buffer[976] = 18'b100000000000000000;
 buffer[977] = 18'b100000000000000000;
 buffer[978] = 18'b100000000000000000;
 buffer[979] = 18'b100000000000000000;
 buffer[980] = 18'b100000000000000000;
 buffer[981] = 18'b100000000000000000;
 buffer[982] = 18'b100000000000000000;
 buffer[983] = 18'b100000000000000000;
 buffer[984] = 18'b100000000000000000;
 buffer[985] = 18'b100000000000000000;
 buffer[986] = 18'b100000000000000000;
 buffer[987] = 18'b100000000000000000;
 buffer[988] = 18'b100000000000000000;
 buffer[989] = 18'b100000000000000000;
 buffer[990] = 18'b100000000000000000;
 buffer[991] = 18'b100000000000000000;
 buffer[992] = 18'b100000000000000000;
 buffer[993] = 18'b100000000000000000;
 buffer[994] = 18'b100000000000000000;
 buffer[995] = 18'b100000000000000000;
 buffer[996] = 18'b100000000000000000;
 buffer[997] = 18'b100000000000000000;
 buffer[998] = 18'b100000000000000000;
 buffer[999] = 18'b100000000000000000;
 buffer[1000] = 18'b100000000000000000;
 buffer[1001] = 18'b100000000000000000;
 buffer[1002] = 18'b100000000000000000;
 buffer[1003] = 18'b100000000000000000;
 buffer[1004] = 18'b100000000000000000;
 buffer[1005] = 18'b100000000000000000;
 buffer[1006] = 18'b100000000000000000;
 buffer[1007] = 18'b100000000000000000;
 buffer[1008] = 18'b100000000000000000;
 buffer[1009] = 18'b100000000000000000;
 buffer[1010] = 18'b100000000000000000;
 buffer[1011] = 18'b100000000000000000;
 buffer[1012] = 18'b100000000000000000;
 buffer[1013] = 18'b100000000000000000;
 buffer[1014] = 18'b100000000000000000;
 buffer[1015] = 18'b100000000000000000;
 buffer[1016] = 18'b100000000000000000;
 buffer[1017] = 18'b100000000000000000;
 buffer[1018] = 18'b100000000000000000;
 buffer[1019] = 18'b100000000000000000;
 buffer[1020] = 18'b100000000000000000;
 buffer[1021] = 18'b100000000000000000;
 buffer[1022] = 18'b100000000000000000;
 buffer[1023] = 18'b100000000000000000;
 buffer[1024] = 18'b100000000000000000;
 buffer[1025] = 18'b100000000000000000;
 buffer[1026] = 18'b100000000000000000;
 buffer[1027] = 18'b100000000000000000;
 buffer[1028] = 18'b100000000000000000;
 buffer[1029] = 18'b100000000000000000;
 buffer[1030] = 18'b100000000000000000;
 buffer[1031] = 18'b100000000000000000;
 buffer[1032] = 18'b100000000000000000;
 buffer[1033] = 18'b100000000000000000;
 buffer[1034] = 18'b100000000000000000;
 buffer[1035] = 18'b100000000000000000;
 buffer[1036] = 18'b100000000000000000;
 buffer[1037] = 18'b100000000000000000;
 buffer[1038] = 18'b100000000000000000;
 buffer[1039] = 18'b100000000000000000;
 buffer[1040] = 18'b100000000000000000;
 buffer[1041] = 18'b100000000000000000;
 buffer[1042] = 18'b100000000000000000;
 buffer[1043] = 18'b100000000000000000;
 buffer[1044] = 18'b100000000000000000;
 buffer[1045] = 18'b100000000000000000;
 buffer[1046] = 18'b100000000000000000;
 buffer[1047] = 18'b100000000000000000;
 buffer[1048] = 18'b100000000000000000;
 buffer[1049] = 18'b100000000000000000;
 buffer[1050] = 18'b100000000000000000;
 buffer[1051] = 18'b100000000000000000;
 buffer[1052] = 18'b100000000000000000;
 buffer[1053] = 18'b100000000000000000;
 buffer[1054] = 18'b100000000000000000;
 buffer[1055] = 18'b100000000000000000;
 buffer[1056] = 18'b100000000000000000;
 buffer[1057] = 18'b100000000000000000;
 buffer[1058] = 18'b100000000000000000;
 buffer[1059] = 18'b100000000000000000;
 buffer[1060] = 18'b100000000000000000;
 buffer[1061] = 18'b100000000000000000;
 buffer[1062] = 18'b100000000000000000;
 buffer[1063] = 18'b100000000000000000;
 buffer[1064] = 18'b100000000000000000;
 buffer[1065] = 18'b100000000000000000;
 buffer[1066] = 18'b100000000000000000;
 buffer[1067] = 18'b100000000000000000;
 buffer[1068] = 18'b100000000000000000;
 buffer[1069] = 18'b100000000000000000;
 buffer[1070] = 18'b100000000000000000;
 buffer[1071] = 18'b100000000000000000;
 buffer[1072] = 18'b100000000000000000;
 buffer[1073] = 18'b100000000000000000;
 buffer[1074] = 18'b100000000000000000;
 buffer[1075] = 18'b100000000000000000;
 buffer[1076] = 18'b100000000000000000;
 buffer[1077] = 18'b100000000000000000;
 buffer[1078] = 18'b100000000000000000;
 buffer[1079] = 18'b100000000000000000;
 buffer[1080] = 18'b100000000000000000;
 buffer[1081] = 18'b100000000000000000;
 buffer[1082] = 18'b100000000000000000;
 buffer[1083] = 18'b100000000000000000;
 buffer[1084] = 18'b100000000000000000;
 buffer[1085] = 18'b100000000000000000;
 buffer[1086] = 18'b100000000000000000;
 buffer[1087] = 18'b100000000000000000;
 buffer[1088] = 18'b100000000000000000;
 buffer[1089] = 18'b100000000000000000;
 buffer[1090] = 18'b100000000000000000;
 buffer[1091] = 18'b100000000000000000;
 buffer[1092] = 18'b100000000000000000;
 buffer[1093] = 18'b100000000000000000;
 buffer[1094] = 18'b100000000000000000;
 buffer[1095] = 18'b100000000000000000;
 buffer[1096] = 18'b100000000000000000;
 buffer[1097] = 18'b100000000000000000;
 buffer[1098] = 18'b100000000000000000;
 buffer[1099] = 18'b100000000000000000;
 buffer[1100] = 18'b100000000000000000;
 buffer[1101] = 18'b100000000000000000;
 buffer[1102] = 18'b100000000000000000;
 buffer[1103] = 18'b100000000000000000;
 buffer[1104] = 18'b100000000000000000;
 buffer[1105] = 18'b100000000000000000;
 buffer[1106] = 18'b100000000000000000;
 buffer[1107] = 18'b100000000000000000;
 buffer[1108] = 18'b100000000000000000;
 buffer[1109] = 18'b100000000000000000;
 buffer[1110] = 18'b100000000000000000;
 buffer[1111] = 18'b100000000000000000;
 buffer[1112] = 18'b100000000000000000;
 buffer[1113] = 18'b100000000000000000;
 buffer[1114] = 18'b100000000000000000;
 buffer[1115] = 18'b100000000000000000;
 buffer[1116] = 18'b100000000000000000;
 buffer[1117] = 18'b100000000000000000;
 buffer[1118] = 18'b100000000000000000;
 buffer[1119] = 18'b100000000000000000;
 buffer[1120] = 18'b100000000000000000;
 buffer[1121] = 18'b100000000000000000;
 buffer[1122] = 18'b100000000000000000;
 buffer[1123] = 18'b100000000000000000;
 buffer[1124] = 18'b100000000000000000;
 buffer[1125] = 18'b100000000000000000;
 buffer[1126] = 18'b100000000000000000;
 buffer[1127] = 18'b100000000000000000;
 buffer[1128] = 18'b100000000000000000;
 buffer[1129] = 18'b100000000000000000;
 buffer[1130] = 18'b100000000000000000;
 buffer[1131] = 18'b100000000000000000;
 buffer[1132] = 18'b100000000000000000;
 buffer[1133] = 18'b100000000000000000;
 buffer[1134] = 18'b100000000000000000;
 buffer[1135] = 18'b100000000000000000;
 buffer[1136] = 18'b100000000000000000;
 buffer[1137] = 18'b100000000000000000;
 buffer[1138] = 18'b100000000000000000;
 buffer[1139] = 18'b100000000000000000;
 buffer[1140] = 18'b100000000000000000;
 buffer[1141] = 18'b100000000000000000;
 buffer[1142] = 18'b100000000000000000;
 buffer[1143] = 18'b100000000000000000;
 buffer[1144] = 18'b100000000000000000;
 buffer[1145] = 18'b100000000000000000;
 buffer[1146] = 18'b100000000000000000;
 buffer[1147] = 18'b100000000000000000;
 buffer[1148] = 18'b100000000000000000;
 buffer[1149] = 18'b100000000000000000;
 buffer[1150] = 18'b100000000000000000;
 buffer[1151] = 18'b100000000000000000;
 buffer[1152] = 18'b100000000000000000;
 buffer[1153] = 18'b100000000000000000;
 buffer[1154] = 18'b100000000000000000;
 buffer[1155] = 18'b100000000000000000;
 buffer[1156] = 18'b100000000000000000;
 buffer[1157] = 18'b100000000000000000;
 buffer[1158] = 18'b100000000000000000;
 buffer[1159] = 18'b100000000000000000;
 buffer[1160] = 18'b100000000000000000;
 buffer[1161] = 18'b100000000000000000;
 buffer[1162] = 18'b100000000000000000;
 buffer[1163] = 18'b100000000000000000;
 buffer[1164] = 18'b100000000000000000;
 buffer[1165] = 18'b100000000000000000;
 buffer[1166] = 18'b100000000000000000;
 buffer[1167] = 18'b100000000000000000;
 buffer[1168] = 18'b100000000000000000;
 buffer[1169] = 18'b100000000000000000;
 buffer[1170] = 18'b100000000000000000;
 buffer[1171] = 18'b100000000000000000;
 buffer[1172] = 18'b100000000000000000;
 buffer[1173] = 18'b100000000000000000;
 buffer[1174] = 18'b100000000000000000;
 buffer[1175] = 18'b100000000000000000;
 buffer[1176] = 18'b100000000000000000;
 buffer[1177] = 18'b100000000000000000;
 buffer[1178] = 18'b100000000000000000;
 buffer[1179] = 18'b100000000000000000;
 buffer[1180] = 18'b100000000000000000;
 buffer[1181] = 18'b100000000000000000;
 buffer[1182] = 18'b100000000000000000;
 buffer[1183] = 18'b100000000000000000;
 buffer[1184] = 18'b100000000000000000;
 buffer[1185] = 18'b100000000000000000;
 buffer[1186] = 18'b100000000000000000;
 buffer[1187] = 18'b100000000000000000;
 buffer[1188] = 18'b100000000000000000;
 buffer[1189] = 18'b100000000000000000;
 buffer[1190] = 18'b100000000000000000;
 buffer[1191] = 18'b100000000000000000;
 buffer[1192] = 18'b100000000000000000;
 buffer[1193] = 18'b100000000000000000;
 buffer[1194] = 18'b100000000000000000;
 buffer[1195] = 18'b100000000000000000;
 buffer[1196] = 18'b100000000000000000;
 buffer[1197] = 18'b100000000000000000;
 buffer[1198] = 18'b100000000000000000;
 buffer[1199] = 18'b100000000000000000;
 buffer[1200] = 18'b100000000000000000;
 buffer[1201] = 18'b100000000000000000;
 buffer[1202] = 18'b100000000000000000;
 buffer[1203] = 18'b100000000000000000;
 buffer[1204] = 18'b100000000000000000;
 buffer[1205] = 18'b100000000000000000;
 buffer[1206] = 18'b100000000000000000;
 buffer[1207] = 18'b100000000000000000;
 buffer[1208] = 18'b100000000000000000;
 buffer[1209] = 18'b100000000000000000;
 buffer[1210] = 18'b100000000000000000;
 buffer[1211] = 18'b100000000000000000;
 buffer[1212] = 18'b100000000000000000;
 buffer[1213] = 18'b100000000000000000;
 buffer[1214] = 18'b100000000000000000;
 buffer[1215] = 18'b100000000000000000;
 buffer[1216] = 18'b100000000000000000;
 buffer[1217] = 18'b100000000000000000;
 buffer[1218] = 18'b100000000000000000;
 buffer[1219] = 18'b100000000000000000;
 buffer[1220] = 18'b100000000000000000;
 buffer[1221] = 18'b100000000000000000;
 buffer[1222] = 18'b100000000000000000;
 buffer[1223] = 18'b100000000000000000;
 buffer[1224] = 18'b100000000000000000;
 buffer[1225] = 18'b100000000000000000;
 buffer[1226] = 18'b100000000000000000;
 buffer[1227] = 18'b100000000000000000;
 buffer[1228] = 18'b100000000000000000;
 buffer[1229] = 18'b100000000000000000;
 buffer[1230] = 18'b100000000000000000;
 buffer[1231] = 18'b100000000000000000;
 buffer[1232] = 18'b100000000000000000;
 buffer[1233] = 18'b100000000000000000;
 buffer[1234] = 18'b100000000000000000;
 buffer[1235] = 18'b100000000000000000;
 buffer[1236] = 18'b100000000000000000;
 buffer[1237] = 18'b100000000000000000;
 buffer[1238] = 18'b100000000000000000;
 buffer[1239] = 18'b100000000000000000;
 buffer[1240] = 18'b100000000000000000;
 buffer[1241] = 18'b100000000000000000;
 buffer[1242] = 18'b100000000000000000;
 buffer[1243] = 18'b100000000000000000;
 buffer[1244] = 18'b100000000000000000;
 buffer[1245] = 18'b100000000000000000;
 buffer[1246] = 18'b100000000000000000;
 buffer[1247] = 18'b100000000000000000;
 buffer[1248] = 18'b100000000000000000;
 buffer[1249] = 18'b100000000000000000;
 buffer[1250] = 18'b100000000000000000;
 buffer[1251] = 18'b100000000000000000;
 buffer[1252] = 18'b100000000000000000;
 buffer[1253] = 18'b100000000000000000;
 buffer[1254] = 18'b100000000000000000;
 buffer[1255] = 18'b100000000000000000;
 buffer[1256] = 18'b100000000000000000;
 buffer[1257] = 18'b100000000000000000;
 buffer[1258] = 18'b100000000000000000;
 buffer[1259] = 18'b100000000000000000;
 buffer[1260] = 18'b100000000000000000;
 buffer[1261] = 18'b100000000000000000;
 buffer[1262] = 18'b100000000000000000;
 buffer[1263] = 18'b100000000000000000;
 buffer[1264] = 18'b100000000000000000;
 buffer[1265] = 18'b100000000000000000;
 buffer[1266] = 18'b100000000000000000;
 buffer[1267] = 18'b100000000000000000;
 buffer[1268] = 18'b100000000000000000;
 buffer[1269] = 18'b100000000000000000;
 buffer[1270] = 18'b100000000000000000;
 buffer[1271] = 18'b100000000000000000;
 buffer[1272] = 18'b100000000000000000;
 buffer[1273] = 18'b100000000000000000;
 buffer[1274] = 18'b100000000000000000;
 buffer[1275] = 18'b100000000000000000;
 buffer[1276] = 18'b100000000000000000;
 buffer[1277] = 18'b100000000000000000;
 buffer[1278] = 18'b100000000000000000;
 buffer[1279] = 18'b100000000000000000;
 buffer[1280] = 18'b100000000000000000;
 buffer[1281] = 18'b100000000000000000;
 buffer[1282] = 18'b100000000000000000;
 buffer[1283] = 18'b100000000000000000;
 buffer[1284] = 18'b100000000000000000;
 buffer[1285] = 18'b100000000000000000;
 buffer[1286] = 18'b100000000000000000;
 buffer[1287] = 18'b100000000000000000;
 buffer[1288] = 18'b100000000000000000;
 buffer[1289] = 18'b100000000000000000;
 buffer[1290] = 18'b100000000000000000;
 buffer[1291] = 18'b100000000000000000;
 buffer[1292] = 18'b100000000000000000;
 buffer[1293] = 18'b100000000000000000;
 buffer[1294] = 18'b100000000000000000;
 buffer[1295] = 18'b100000000000000000;
 buffer[1296] = 18'b100000000000000000;
 buffer[1297] = 18'b100000000000000000;
 buffer[1298] = 18'b100000000000000000;
 buffer[1299] = 18'b100000000000000000;
 buffer[1300] = 18'b100000000000000000;
 buffer[1301] = 18'b100000000000000000;
 buffer[1302] = 18'b100000000000000000;
 buffer[1303] = 18'b100000000000000000;
 buffer[1304] = 18'b100000000000000000;
 buffer[1305] = 18'b100000000000000000;
 buffer[1306] = 18'b100000000000000000;
 buffer[1307] = 18'b100000000000000000;
 buffer[1308] = 18'b100000000000000000;
 buffer[1309] = 18'b100000000000000000;
 buffer[1310] = 18'b100000000000000000;
 buffer[1311] = 18'b100000000000000000;
 buffer[1312] = 18'b100000000000000000;
 buffer[1313] = 18'b100000000000000000;
 buffer[1314] = 18'b100000000000000000;
 buffer[1315] = 18'b100000000000000000;
 buffer[1316] = 18'b100000000000000000;
 buffer[1317] = 18'b100000000000000000;
 buffer[1318] = 18'b100000000000000000;
 buffer[1319] = 18'b100000000000000000;
 buffer[1320] = 18'b100000000000000000;
 buffer[1321] = 18'b100000000000000000;
 buffer[1322] = 18'b100000000000000000;
 buffer[1323] = 18'b100000000000000000;
 buffer[1324] = 18'b100000000000000000;
 buffer[1325] = 18'b100000000000000000;
 buffer[1326] = 18'b100000000000000000;
 buffer[1327] = 18'b100000000000000000;
 buffer[1328] = 18'b100000000000000000;
 buffer[1329] = 18'b100000000000000000;
 buffer[1330] = 18'b100000000000000000;
 buffer[1331] = 18'b100000000000000000;
 buffer[1332] = 18'b100000000000000000;
 buffer[1333] = 18'b100000000000000000;
 buffer[1334] = 18'b100000000000000000;
 buffer[1335] = 18'b100000000000000000;
 buffer[1336] = 18'b100000000000000000;
 buffer[1337] = 18'b100000000000000000;
 buffer[1338] = 18'b100000000000000000;
 buffer[1339] = 18'b100000000000000000;
 buffer[1340] = 18'b100000000000000000;
 buffer[1341] = 18'b100000000000000000;
 buffer[1342] = 18'b100000000000000000;
 buffer[1343] = 18'b100000000000000000;
end

endmodule

module M_tilemap (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_tm_x,
in_tm_y,
in_tm_character,
in_tm_foreground,
in_tm_background,
in_tm_write,
in_tile_writer_tile,
in_tile_writer_line,
in_tile_writer_bitmap,
in_tm_scrollwrap,
out_pix_red,
out_pix_green,
out_pix_blue,
out_tilemap_display,
out_tm_lastaction,
out_tm_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [5:0] in_tm_x;
input  [5:0] in_tm_y;
input  [4:0] in_tm_character;
input  [5:0] in_tm_foreground;
input  [6:0] in_tm_background;
input  [0:0] in_tm_write;
input  [4:0] in_tile_writer_tile;
input  [3:0] in_tile_writer_line;
input  [15:0] in_tile_writer_bitmap;
input  [3:0] in_tm_scrollwrap;
output  [1:0] out_pix_red;
output  [1:0] out_pix_green;
output  [1:0] out_pix_blue;
output  [0:0] out_tilemap_display;
output  [3:0] out_tm_lastaction;
output  [1:0] out_tm_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [15:0] _w_mem_tiles16x16_rdata0;
wire  [17:0] _w_mem_tiles_rdata0;
wire  [17:0] _w_mem_tiles_copy_rdata0;
reg  [10:0] _t_tiles_addr0;
reg  [0:0] _t_tiles_wenable1;
reg  [17:0] _t_tiles_wdata1;
reg  [10:0] _t_tiles_addr1;
reg  [10:0] _t_tiles_copy_addr0;
reg  [0:0] _t_tiles_copy_wenable1;
reg  [17:0] _t_tiles_copy_wdata1;
reg  [10:0] _t_tiles_copy_addr1;
wire  [10:0] _w_xtmpos;
wire  [10:0] _w_ytmpos;
wire  [3:0] _w_xintm;
wire  [3:0] _w_yintm;
wire  [0:0] _w_tmpixel;

reg  [8:0] _d_tiles16x16_addr0;
reg  [8:0] _q_tiles16x16_addr0;
reg  [0:0] _d_tiles16x16_wenable1;
reg  [0:0] _q_tiles16x16_wenable1;
reg  [15:0] _d_tiles16x16_wdata1;
reg  [15:0] _q_tiles16x16_wdata1;
reg  [8:0] _d_tiles16x16_addr1;
reg  [8:0] _q_tiles16x16_addr1;
reg signed [4:0] _d_tm_offset_x;
reg signed [4:0] _q_tm_offset_x;
reg signed [4:0] _d_tm_offset_y;
reg signed [4:0] _q_tm_offset_y;
reg  [0:0] _d_tm_scroll;
reg  [0:0] _q_tm_scroll;
reg  [0:0] _d_tm_goleft;
reg  [0:0] _q_tm_goleft;
reg  [0:0] _d_tm_goup;
reg  [0:0] _q_tm_goup;
reg  [5:0] _d_x_cursor;
reg  [5:0] _q_x_cursor;
reg  [5:0] _d_y_cursor;
reg  [5:0] _q_y_cursor;
reg  [10:0] _d_y_cursor_addr;
reg  [10:0] _q_y_cursor_addr;
reg  [17:0] _d_new_tile;
reg  [17:0] _q_new_tile;
reg  [10:0] _d_tmcsaddr;
reg  [10:0] _q_tmcsaddr;
reg  [1:0] _d_pix_red,_q_pix_red;
reg  [1:0] _d_pix_green,_q_pix_green;
reg  [1:0] _d_pix_blue,_q_pix_blue;
reg  [0:0] _d_tilemap_display,_q_tilemap_display;
reg  [3:0] _d_tm_lastaction,_q_tm_lastaction;
reg  [1:0] _d_tm_active,_q_tm_active;
reg  [4:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_tilemap_display = _d_tilemap_display;
assign out_tm_lastaction = _q_tm_lastaction;
assign out_tm_active = _q_tm_active;
assign out_done = (_q_index == 22);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_tiles16x16_addr0 <= 0;
_q_tiles16x16_wenable1 <= 0;
_q_tiles16x16_wdata1 <= 0;
_q_tiles16x16_addr1 <= 0;
_q_tm_offset_x <= 0;
_q_tm_offset_y <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_tiles16x16_addr0 <= _d_tiles16x16_addr0;
_q_tiles16x16_wenable1 <= _d_tiles16x16_wenable1;
_q_tiles16x16_wdata1 <= _d_tiles16x16_wdata1;
_q_tiles16x16_addr1 <= _d_tiles16x16_addr1;
_q_tm_offset_x <= _d_tm_offset_x;
_q_tm_offset_y <= _d_tm_offset_y;
_q_tm_scroll <= _d_tm_scroll;
_q_tm_goleft <= _d_tm_goleft;
_q_tm_goup <= _d_tm_goup;
_q_x_cursor <= _d_x_cursor;
_q_y_cursor <= _d_y_cursor;
_q_y_cursor_addr <= _d_y_cursor_addr;
_q_new_tile <= _d_new_tile;
_q_tmcsaddr <= _d_tmcsaddr;
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_tilemap_display <= _d_tilemap_display;
_q_tm_lastaction <= _d_tm_lastaction;
_q_tm_active <= _d_tm_active;
_q_index <= _d_index;
  end
end


M_tilemap_mem_tiles16x16 __mem__tiles16x16(
.clock0(clock),
.clock1(clock),
.in_tiles16x16_addr0(_d_tiles16x16_addr0),
.in_tiles16x16_wenable1(_d_tiles16x16_wenable1),
.in_tiles16x16_wdata1(_d_tiles16x16_wdata1),
.in_tiles16x16_addr1(_d_tiles16x16_addr1),
.out_tiles16x16_rdata0(_w_mem_tiles16x16_rdata0)
);
M_tilemap_mem_tiles __mem__tiles(
.clock0(clock),
.clock1(clock),
.in_tiles_addr0(_t_tiles_addr0),
.in_tiles_wenable1(_t_tiles_wenable1),
.in_tiles_wdata1(_t_tiles_wdata1),
.in_tiles_addr1(_t_tiles_addr1),
.out_tiles_rdata0(_w_mem_tiles_rdata0)
);
M_tilemap_mem_tiles_copy __mem__tiles_copy(
.clock0(clock),
.clock1(clock),
.in_tiles_copy_addr0(_t_tiles_copy_addr0),
.in_tiles_copy_wenable1(_t_tiles_copy_wenable1),
.in_tiles_copy_wdata1(_t_tiles_copy_wdata1),
.in_tiles_copy_addr1(_t_tiles_copy_addr1),
.out_tiles_copy_rdata0(_w_mem_tiles_copy_rdata0)
);

assign _w_tmpixel = _w_mem_tiles16x16_rdata0[15-_w_xintm+:1];
assign _w_yintm = {1'b0,(in_pix_y)&15}+_d_tm_offset_y;
assign _w_xintm = {1'b0,(in_pix_x)&15}+_d_tm_offset_x;
assign _w_ytmpos = ((in_pix_vblank?(11'd16+{{6{_d_tm_offset_y[4+:1]}},_d_tm_offset_y}):in_pix_y+(11'd16+{{6{_d_tm_offset_y[4+:1]}},_d_tm_offset_y}))>>4)*42;
assign _w_xtmpos = (in_pix_active?in_pix_x+(11'd18+{{6{_d_tm_offset_x[4+:1]}},_d_tm_offset_x}):(11'd16+{{6{_d_tm_offset_x[4+:1]}},_d_tm_offset_x}))>>4;

always @* begin
_d_tiles16x16_addr0 = _q_tiles16x16_addr0;
_d_tiles16x16_wenable1 = _q_tiles16x16_wenable1;
_d_tiles16x16_wdata1 = _q_tiles16x16_wdata1;
_d_tiles16x16_addr1 = _q_tiles16x16_addr1;
_d_tm_offset_x = _q_tm_offset_x;
_d_tm_offset_y = _q_tm_offset_y;
_d_tm_scroll = _q_tm_scroll;
_d_tm_goleft = _q_tm_goleft;
_d_tm_goup = _q_tm_goup;
_d_x_cursor = _q_x_cursor;
_d_y_cursor = _q_y_cursor;
_d_y_cursor_addr = _q_y_cursor_addr;
_d_new_tile = _q_new_tile;
_d_tmcsaddr = _q_tmcsaddr;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_tilemap_display = _q_tilemap_display;
_d_tm_lastaction = _q_tm_lastaction;
_d_tm_active = _q_tm_active;
_d_index = _q_index;
_t_tiles_addr0 = 0;
_t_tiles_wenable1 = 0;
_t_tiles_wdata1 = 0;
_t_tiles_addr1 = 0;
_t_tiles_copy_addr0 = 0;
_t_tiles_copy_wenable1 = 0;
_t_tiles_copy_wdata1 = 0;
_t_tiles_copy_addr1 = 0;
// _always_pre
_t_tiles_addr0 = _w_xtmpos+_w_ytmpos;
_t_tiles_wenable1 = 1;
_t_tiles_copy_wenable1 = 1;
_d_tiles16x16_addr0 = _w_mem_tiles_rdata0[0+:5]*16+_w_yintm;
_d_tiles16x16_addr1 = in_tile_writer_tile*16+in_tile_writer_line;
_d_tiles16x16_wdata1 = in_tile_writer_bitmap;
_d_tiles16x16_wenable1 = 1;
_d_tilemap_display = in_pix_active&&((_w_tmpixel)||(~_w_mem_tiles_rdata0[17+:1]));
_d_pix_red = _w_tmpixel?_w_mem_tiles_rdata0[9+:2]:_w_mem_tiles_rdata0[15+:2];
_d_pix_green = _w_tmpixel?_w_mem_tiles_rdata0[7+:2]:_w_mem_tiles_rdata0[13+:2];
_d_pix_blue = _w_tmpixel?_w_mem_tiles_rdata0[5+:2]:_w_mem_tiles_rdata0[11+:2];
_d_index = 22;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_tiles16x16_addr0 = 0;
_d_tiles16x16_wenable1 = 0;
_d_tiles16x16_wdata1 = 0;
_d_tiles16x16_addr1 = 0;
_t_tiles_addr0 = 0;
_t_tiles_wenable1 = 0;
_t_tiles_wdata1 = 0;
_t_tiles_addr1 = 0;
_t_tiles_copy_addr0 = 0;
_t_tiles_copy_wenable1 = 0;
_t_tiles_copy_wdata1 = 0;
_t_tiles_copy_addr1 = 0;
_d_tm_offset_x = 0;
_d_tm_offset_y = 0;
// --
_t_tiles_addr1 = 0;
_t_tiles_wdata1 = {1'b1,6'b0,6'b0,5'b0};
_t_tiles_copy_addr1 = 0;
_t_tiles_copy_wdata1 = {1'b1,6'b0,6'b0,5'b0};
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_tm_write==1) begin
// __block_5
// __block_7
_t_tiles_addr1 = in_tm_x+in_tm_y*42;
_t_tiles_wdata1 = {in_tm_background,in_tm_foreground,in_tm_character};
_t_tiles_copy_addr1 = in_tm_x+in_tm_y*42;
_t_tiles_copy_wdata1 = {in_tm_background,in_tm_foreground,in_tm_character};
// __block_8
end else begin
// __block_6
end
// __block_9
  case (_q_tm_active)
  0: begin
// __block_11_case
// __block_12
  case (in_tm_scrollwrap)
  1: begin
// __block_14_case
// __block_15
if (_q_tm_offset_x==15) begin
// __block_16
// __block_18
_d_tm_scroll = 1;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goleft = 1;
_d_tm_active = 1;
// __block_19
end else begin
// __block_17
// __block_20
_d_tm_offset_x = _q_tm_offset_x+1;
_d_tm_lastaction = 0;
// __block_21
end
// __block_22
// __block_23
  end
  2: begin
// __block_24_case
// __block_25
if (_q_tm_offset_y==15) begin
// __block_26
// __block_28
_d_tm_scroll = 1;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goup = 1;
_d_tm_active = 2;
// __block_29
end else begin
// __block_27
// __block_30
_d_tm_offset_y = _q_tm_offset_y+1;
_d_tm_lastaction = 0;
// __block_31
end
// __block_32
// __block_33
  end
  3: begin
// __block_34_case
// __block_35
if (_q_tm_offset_x==-15) begin
// __block_36
// __block_38
_d_tm_scroll = 1;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goleft = 0;
_d_tm_active = 1;
// __block_39
end else begin
// __block_37
// __block_40
_d_tm_offset_x = _q_tm_offset_x-1;
_d_tm_lastaction = 0;
// __block_41
end
// __block_42
// __block_43
  end
  4: begin
// __block_44_case
// __block_45
if (_q_tm_offset_y==-15) begin
// __block_46
// __block_48
_d_tm_scroll = 1;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goup = 0;
_d_tm_active = 2;
// __block_49
end else begin
// __block_47
// __block_50
_d_tm_offset_y = _q_tm_offset_y-1;
_d_tm_lastaction = 0;
// __block_51
end
// __block_52
// __block_53
  end
  5: begin
// __block_54_case
// __block_55
if (_q_tm_offset_x==15) begin
// __block_56
// __block_58
_d_tm_scroll = 0;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goleft = 1;
_d_tm_active = 1;
// __block_59
end else begin
// __block_57
// __block_60
_d_tm_offset_x = _q_tm_offset_x+1;
_d_tm_lastaction = 0;
// __block_61
end
// __block_62
// __block_63
  end
  6: begin
// __block_64_case
// __block_65
if (_q_tm_offset_y==15) begin
// __block_66
// __block_68
_d_tm_scroll = 0;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goup = 1;
_d_tm_active = 2;
// __block_69
end else begin
// __block_67
// __block_70
_d_tm_offset_y = _q_tm_offset_y+1;
_d_tm_lastaction = 0;
// __block_71
end
// __block_72
// __block_73
  end
  7: begin
// __block_74_case
// __block_75
if (_q_tm_offset_x==-15) begin
// __block_76
// __block_78
_d_tm_scroll = 0;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goleft = 0;
_d_tm_active = 1;
// __block_79
end else begin
// __block_77
// __block_80
_d_tm_offset_x = _q_tm_offset_x-1;
_d_tm_lastaction = 0;
// __block_81
end
// __block_82
// __block_83
  end
  8: begin
// __block_84_case
// __block_85
if (_q_tm_offset_y==-15) begin
// __block_86
// __block_88
_d_tm_scroll = 0;
_d_tm_lastaction = in_tm_scrollwrap;
_d_tm_goup = 0;
_d_tm_active = 2;
// __block_89
end else begin
// __block_87
// __block_90
_d_tm_offset_y = _q_tm_offset_y-1;
_d_tm_lastaction = 0;
// __block_91
end
// __block_92
// __block_93
  end
  9: begin
// __block_94_case
// __block_95
_d_tm_active = 3;
_d_tm_lastaction = 9;
// __block_96
  end
endcase
// __block_13
// __block_97
_d_index = 1;
  end
  1: begin
// __block_98_case
// __block_99
_d_y_cursor = 0;
_d_y_cursor_addr = 0;
_d_index = 3;
  end
  2: begin
// __block_117_case
// __block_118
_d_x_cursor = 0;
_d_index = 4;
  end
  3: begin
// __block_135_case
// __block_136
_d_tmcsaddr = 0;
_d_index = 5;
  end
endcase
end else begin
_d_index = 2;
end
end
3: begin
// __block_100
_d_index = 6;
end
4: begin
// __block_119
_d_index = 7;
end
5: begin
// __block_137
_d_index = 8;
end
2: begin
// __block_3
_d_index = 22;
end
6: begin
// __while__block_101
if (_q_y_cursor<32) begin
// __block_102
// __block_104
_d_x_cursor = _q_tm_goleft?0:41;
_t_tiles_copy_addr0 = _q_tm_goleft?_q_y_cursor_addr:41+_q_y_cursor_addr;
_d_index = 12;
end else begin
_d_index = 9;
end
end
7: begin
// __while__block_120
if (_q_x_cursor<42) begin
// __block_121
// __block_123
_d_y_cursor = _q_tm_goup?0:31;
_d_y_cursor_addr = _q_tm_goup?0:1302;
_t_tiles_copy_addr0 = _q_x_cursor;
_d_index = 13;
end else begin
_d_index = 10;
end
end
8: begin
// __while__block_138
if (_q_tmcsaddr<1344) begin
// __block_139
// __block_141
_t_tiles_addr1 = _q_tmcsaddr;
_t_tiles_wdata1 = {1'b1,6'b0,6'b0,5'b0};
_t_tiles_copy_addr1 = _q_tmcsaddr;
_t_tiles_copy_wdata1 = {1'b1,6'b0,6'b0,5'b0};
_d_tmcsaddr = _q_tmcsaddr+1;
// __block_142
_d_index = 8;
end else begin
_d_index = 11;
end
end
12: begin
// __block_105
_d_new_tile = (_q_tm_scroll==1)?{1'b1,6'b0,6'b0,5'b0}:_w_mem_tiles_copy_rdata0;
_d_index = 14;
end
9: begin
// __block_115
_d_tm_offset_x = 0;
_d_tm_active = 0;
// __block_116
_d_index = 1;
end
13: begin
// __block_124
_d_new_tile = (_q_tm_scroll==1)?{1'b1,6'b0,6'b0,5'b0}:_w_mem_tiles_copy_rdata0;
_d_index = 15;
end
10: begin
// __block_133
_d_tm_offset_y = 0;
_d_tm_active = 0;
// __block_134
_d_index = 1;
end
11: begin
// __block_143
_d_tm_offset_x = 0;
_d_tm_offset_y = 0;
_d_tm_active = 0;
// __block_144
_d_index = 1;
end
14: begin
// __block_106
_d_index = 16;
end
15: begin
// __block_125
_d_index = 17;
end
16: begin
// __while__block_107
if (_q_tm_goleft?(_q_x_cursor<42):(_q_x_cursor>0)) begin
// __block_108
// __block_110
_t_tiles_copy_addr0 = _q_tm_goleft?(_q_x_cursor+1+_q_y_cursor_addr):(_q_x_cursor-1+_q_y_cursor_addr);
_d_index = 20;
end else begin
_d_index = 18;
end
end
17: begin
// __while__block_126
if (_q_tm_goup?(_q_y_cursor<31):(_q_y_cursor>0)) begin
// __block_127
// __block_129
_t_tiles_copy_addr0 = _q_tm_goup?(_q_x_cursor+_q_y_cursor_addr+42):(_q_x_cursor+_q_y_cursor_addr-42);
_d_index = 21;
end else begin
_d_index = 19;
end
end
20: begin
// __block_111
_t_tiles_addr1 = _q_x_cursor+_q_y_cursor_addr;
_t_tiles_wdata1 = _w_mem_tiles_copy_rdata0;
_t_tiles_copy_addr1 = _q_x_cursor+_q_y_cursor_addr;
_t_tiles_copy_wdata1 = _w_mem_tiles_copy_rdata0;
_d_x_cursor = _q_tm_goleft?(_q_x_cursor+1):(_q_x_cursor-1);
// __block_112
_d_index = 16;
end
18: begin
// __block_113
_t_tiles_addr1 = _q_tm_goleft?(41+_q_y_cursor_addr):(_q_y_cursor_addr);
_t_tiles_wdata1 = _q_new_tile;
_t_tiles_copy_addr1 = _q_tm_goleft?(41+_q_y_cursor_addr):(_q_y_cursor_addr);
_t_tiles_copy_wdata1 = _q_new_tile;
_d_y_cursor = _q_y_cursor+1;
_d_y_cursor_addr = _q_y_cursor_addr+42;
// __block_114
_d_index = 6;
end
21: begin
// __block_130
_t_tiles_addr1 = _q_x_cursor+_q_y_cursor_addr;
_t_tiles_wdata1 = _w_mem_tiles_copy_rdata0;
_t_tiles_copy_addr1 = _q_x_cursor+_q_y_cursor_addr;
_t_tiles_copy_wdata1 = _w_mem_tiles_copy_rdata0;
_d_y_cursor = _q_tm_goup?(_q_y_cursor+1):(_q_y_cursor-1);
_d_y_cursor_addr = _q_tm_goup?(_q_y_cursor_addr+42):(_q_y_cursor_addr-42);
// __block_131
_d_index = 17;
end
19: begin
// __block_128
_t_tiles_addr1 = _q_tm_goup?(_q_x_cursor+1302):(_q_x_cursor);
_t_tiles_wdata1 = _q_new_tile;
_t_tiles_copy_addr1 = _q_tm_goup?(_q_x_cursor+1302):(_q_x_cursor);
_t_tiles_copy_wdata1 = _q_new_tile;
_d_x_cursor = _q_x_cursor+1;
// __block_132
_d_index = 7;
end
22: begin // end of tilemap
end
default: begin 
_d_index = 22;
 end
endcase
end
endmodule


module M_apu_mem_waveformtable_1(
input                  [8:0] in_waveformtable_1_addr,
output reg  [3:0] out_waveformtable_1_rdata,
input                                   clock
);
reg  [3:0] buffer[511:0];
always @(posedge clock) begin
   out_waveformtable_1_rdata <= buffer[in_waveformtable_1_addr];
end
initial begin
 buffer[0] = 15;
 buffer[1] = 15;
 buffer[2] = 15;
 buffer[3] = 15;
 buffer[4] = 15;
 buffer[5] = 15;
 buffer[6] = 15;
 buffer[7] = 15;
 buffer[8] = 15;
 buffer[9] = 15;
 buffer[10] = 15;
 buffer[11] = 15;
 buffer[12] = 15;
 buffer[13] = 15;
 buffer[14] = 15;
 buffer[15] = 15;
 buffer[16] = 0;
 buffer[17] = 0;
 buffer[18] = 0;
 buffer[19] = 0;
 buffer[20] = 0;
 buffer[21] = 0;
 buffer[22] = 0;
 buffer[23] = 0;
 buffer[24] = 0;
 buffer[25] = 0;
 buffer[26] = 0;
 buffer[27] = 0;
 buffer[28] = 0;
 buffer[29] = 0;
 buffer[30] = 0;
 buffer[31] = 0;
 buffer[32] = 0;
 buffer[33] = 0;
 buffer[34] = 1;
 buffer[35] = 1;
 buffer[36] = 2;
 buffer[37] = 2;
 buffer[38] = 3;
 buffer[39] = 3;
 buffer[40] = 4;
 buffer[41] = 4;
 buffer[42] = 5;
 buffer[43] = 5;
 buffer[44] = 6;
 buffer[45] = 6;
 buffer[46] = 7;
 buffer[47] = 7;
 buffer[48] = 8;
 buffer[49] = 8;
 buffer[50] = 9;
 buffer[51] = 9;
 buffer[52] = 10;
 buffer[53] = 10;
 buffer[54] = 11;
 buffer[55] = 11;
 buffer[56] = 12;
 buffer[57] = 12;
 buffer[58] = 13;
 buffer[59] = 13;
 buffer[60] = 14;
 buffer[61] = 14;
 buffer[62] = 15;
 buffer[63] = 15;
 buffer[64] = 0;
 buffer[65] = 1;
 buffer[66] = 2;
 buffer[67] = 3;
 buffer[68] = 4;
 buffer[69] = 5;
 buffer[70] = 6;
 buffer[71] = 7;
 buffer[72] = 8;
 buffer[73] = 9;
 buffer[74] = 10;
 buffer[75] = 11;
 buffer[76] = 12;
 buffer[77] = 13;
 buffer[78] = 14;
 buffer[79] = 15;
 buffer[80] = 15;
 buffer[81] = 14;
 buffer[82] = 13;
 buffer[83] = 12;
 buffer[84] = 11;
 buffer[85] = 10;
 buffer[86] = 9;
 buffer[87] = 8;
 buffer[88] = 7;
 buffer[89] = 6;
 buffer[90] = 5;
 buffer[91] = 4;
 buffer[92] = 3;
 buffer[93] = 2;
 buffer[94] = 1;
 buffer[95] = 0;
 buffer[96] = 7;
 buffer[97] = 8;
 buffer[98] = 10;
 buffer[99] = 11;
 buffer[100] = 12;
 buffer[101] = 13;
 buffer[102] = 13;
 buffer[103] = 14;
 buffer[104] = 15;
 buffer[105] = 14;
 buffer[106] = 13;
 buffer[107] = 13;
 buffer[108] = 12;
 buffer[109] = 11;
 buffer[110] = 10;
 buffer[111] = 8;
 buffer[112] = 7;
 buffer[113] = 6;
 buffer[114] = 4;
 buffer[115] = 3;
 buffer[116] = 2;
 buffer[117] = 1;
 buffer[118] = 1;
 buffer[119] = 0;
 buffer[120] = 0;
 buffer[121] = 0;
 buffer[122] = 1;
 buffer[123] = 1;
 buffer[124] = 2;
 buffer[125] = 3;
 buffer[126] = 4;
 buffer[127] = 6;
 buffer[128] = 1;
 buffer[129] = 1;
 buffer[130] = 1;
 buffer[131] = 1;
 buffer[132] = 1;
 buffer[133] = 1;
 buffer[134] = 1;
 buffer[135] = 1;
 buffer[136] = 1;
 buffer[137] = 1;
 buffer[138] = 1;
 buffer[139] = 1;
 buffer[140] = 1;
 buffer[141] = 1;
 buffer[142] = 1;
 buffer[143] = 1;
 buffer[144] = 1;
 buffer[145] = 1;
 buffer[146] = 1;
 buffer[147] = 1;
 buffer[148] = 1;
 buffer[149] = 1;
 buffer[150] = 1;
 buffer[151] = 1;
 buffer[152] = 1;
 buffer[153] = 1;
 buffer[154] = 1;
 buffer[155] = 1;
 buffer[156] = 1;
 buffer[157] = 1;
 buffer[158] = 1;
 buffer[159] = 1;
 buffer[160] = 1;
 buffer[161] = 1;
 buffer[162] = 1;
 buffer[163] = 1;
 buffer[164] = 1;
 buffer[165] = 1;
 buffer[166] = 1;
 buffer[167] = 1;
 buffer[168] = 1;
 buffer[169] = 1;
 buffer[170] = 1;
 buffer[171] = 1;
 buffer[172] = 1;
 buffer[173] = 1;
 buffer[174] = 1;
 buffer[175] = 1;
 buffer[176] = 1;
 buffer[177] = 1;
 buffer[178] = 1;
 buffer[179] = 1;
 buffer[180] = 1;
 buffer[181] = 1;
 buffer[182] = 1;
 buffer[183] = 1;
 buffer[184] = 1;
 buffer[185] = 1;
 buffer[186] = 1;
 buffer[187] = 1;
 buffer[188] = 1;
 buffer[189] = 1;
 buffer[190] = 1;
 buffer[191] = 1;
 buffer[192] = 1;
 buffer[193] = 1;
 buffer[194] = 1;
 buffer[195] = 1;
 buffer[196] = 1;
 buffer[197] = 1;
 buffer[198] = 1;
 buffer[199] = 1;
 buffer[200] = 1;
 buffer[201] = 1;
 buffer[202] = 1;
 buffer[203] = 1;
 buffer[204] = 1;
 buffer[205] = 1;
 buffer[206] = 1;
 buffer[207] = 1;
 buffer[208] = 1;
 buffer[209] = 1;
 buffer[210] = 1;
 buffer[211] = 1;
 buffer[212] = 1;
 buffer[213] = 1;
 buffer[214] = 1;
 buffer[215] = 1;
 buffer[216] = 1;
 buffer[217] = 1;
 buffer[218] = 1;
 buffer[219] = 1;
 buffer[220] = 1;
 buffer[221] = 1;
 buffer[222] = 1;
 buffer[223] = 1;
 buffer[224] = 1;
 buffer[225] = 1;
 buffer[226] = 1;
 buffer[227] = 1;
 buffer[228] = 1;
 buffer[229] = 1;
 buffer[230] = 1;
 buffer[231] = 1;
 buffer[232] = 1;
 buffer[233] = 1;
 buffer[234] = 1;
 buffer[235] = 1;
 buffer[236] = 1;
 buffer[237] = 1;
 buffer[238] = 1;
 buffer[239] = 1;
 buffer[240] = 1;
 buffer[241] = 1;
 buffer[242] = 1;
 buffer[243] = 1;
 buffer[244] = 1;
 buffer[245] = 1;
 buffer[246] = 1;
 buffer[247] = 1;
 buffer[248] = 1;
 buffer[249] = 1;
 buffer[250] = 1;
 buffer[251] = 1;
 buffer[252] = 1;
 buffer[253] = 1;
 buffer[254] = 1;
 buffer[255] = 1;
 buffer[256] = 1;
 buffer[257] = 1;
 buffer[258] = 1;
 buffer[259] = 1;
 buffer[260] = 1;
 buffer[261] = 1;
 buffer[262] = 1;
 buffer[263] = 1;
 buffer[264] = 1;
 buffer[265] = 1;
 buffer[266] = 1;
 buffer[267] = 1;
 buffer[268] = 1;
 buffer[269] = 1;
 buffer[270] = 1;
 buffer[271] = 1;
 buffer[272] = 1;
 buffer[273] = 1;
 buffer[274] = 1;
 buffer[275] = 1;
 buffer[276] = 1;
 buffer[277] = 1;
 buffer[278] = 1;
 buffer[279] = 1;
 buffer[280] = 1;
 buffer[281] = 1;
 buffer[282] = 1;
 buffer[283] = 1;
 buffer[284] = 1;
 buffer[285] = 1;
 buffer[286] = 1;
 buffer[287] = 1;
 buffer[288] = 1;
 buffer[289] = 1;
 buffer[290] = 1;
 buffer[291] = 1;
 buffer[292] = 1;
 buffer[293] = 1;
 buffer[294] = 1;
 buffer[295] = 1;
 buffer[296] = 1;
 buffer[297] = 1;
 buffer[298] = 1;
 buffer[299] = 1;
 buffer[300] = 1;
 buffer[301] = 1;
 buffer[302] = 1;
 buffer[303] = 1;
 buffer[304] = 1;
 buffer[305] = 1;
 buffer[306] = 1;
 buffer[307] = 1;
 buffer[308] = 1;
 buffer[309] = 1;
 buffer[310] = 1;
 buffer[311] = 1;
 buffer[312] = 1;
 buffer[313] = 1;
 buffer[314] = 1;
 buffer[315] = 1;
 buffer[316] = 1;
 buffer[317] = 1;
 buffer[318] = 1;
 buffer[319] = 1;
 buffer[320] = 1;
 buffer[321] = 1;
 buffer[322] = 1;
 buffer[323] = 1;
 buffer[324] = 1;
 buffer[325] = 1;
 buffer[326] = 1;
 buffer[327] = 1;
 buffer[328] = 1;
 buffer[329] = 1;
 buffer[330] = 1;
 buffer[331] = 1;
 buffer[332] = 1;
 buffer[333] = 1;
 buffer[334] = 1;
 buffer[335] = 1;
 buffer[336] = 1;
 buffer[337] = 1;
 buffer[338] = 1;
 buffer[339] = 1;
 buffer[340] = 1;
 buffer[341] = 1;
 buffer[342] = 1;
 buffer[343] = 1;
 buffer[344] = 1;
 buffer[345] = 1;
 buffer[346] = 1;
 buffer[347] = 1;
 buffer[348] = 1;
 buffer[349] = 1;
 buffer[350] = 1;
 buffer[351] = 1;
 buffer[352] = 1;
 buffer[353] = 1;
 buffer[354] = 1;
 buffer[355] = 1;
 buffer[356] = 1;
 buffer[357] = 1;
 buffer[358] = 1;
 buffer[359] = 1;
 buffer[360] = 1;
 buffer[361] = 1;
 buffer[362] = 1;
 buffer[363] = 1;
 buffer[364] = 1;
 buffer[365] = 1;
 buffer[366] = 1;
 buffer[367] = 1;
 buffer[368] = 1;
 buffer[369] = 1;
 buffer[370] = 1;
 buffer[371] = 1;
 buffer[372] = 1;
 buffer[373] = 1;
 buffer[374] = 1;
 buffer[375] = 1;
 buffer[376] = 1;
 buffer[377] = 1;
 buffer[378] = 1;
 buffer[379] = 1;
 buffer[380] = 1;
 buffer[381] = 1;
 buffer[382] = 1;
 buffer[383] = 1;
 buffer[384] = 1;
 buffer[385] = 1;
 buffer[386] = 1;
 buffer[387] = 1;
 buffer[388] = 1;
 buffer[389] = 1;
 buffer[390] = 1;
 buffer[391] = 1;
 buffer[392] = 1;
 buffer[393] = 1;
 buffer[394] = 1;
 buffer[395] = 1;
 buffer[396] = 1;
 buffer[397] = 1;
 buffer[398] = 1;
 buffer[399] = 1;
 buffer[400] = 1;
 buffer[401] = 1;
 buffer[402] = 1;
 buffer[403] = 1;
 buffer[404] = 1;
 buffer[405] = 1;
 buffer[406] = 1;
 buffer[407] = 1;
 buffer[408] = 1;
 buffer[409] = 1;
 buffer[410] = 1;
 buffer[411] = 1;
 buffer[412] = 1;
 buffer[413] = 1;
 buffer[414] = 1;
 buffer[415] = 1;
 buffer[416] = 1;
 buffer[417] = 1;
 buffer[418] = 1;
 buffer[419] = 1;
 buffer[420] = 1;
 buffer[421] = 1;
 buffer[422] = 1;
 buffer[423] = 1;
 buffer[424] = 1;
 buffer[425] = 1;
 buffer[426] = 1;
 buffer[427] = 1;
 buffer[428] = 1;
 buffer[429] = 1;
 buffer[430] = 1;
 buffer[431] = 1;
 buffer[432] = 1;
 buffer[433] = 1;
 buffer[434] = 1;
 buffer[435] = 1;
 buffer[436] = 1;
 buffer[437] = 1;
 buffer[438] = 1;
 buffer[439] = 1;
 buffer[440] = 1;
 buffer[441] = 1;
 buffer[442] = 1;
 buffer[443] = 1;
 buffer[444] = 1;
 buffer[445] = 1;
 buffer[446] = 1;
 buffer[447] = 1;
 buffer[448] = 1;
 buffer[449] = 1;
 buffer[450] = 1;
 buffer[451] = 1;
 buffer[452] = 1;
 buffer[453] = 1;
 buffer[454] = 1;
 buffer[455] = 1;
 buffer[456] = 1;
 buffer[457] = 1;
 buffer[458] = 1;
 buffer[459] = 1;
 buffer[460] = 1;
 buffer[461] = 1;
 buffer[462] = 1;
 buffer[463] = 1;
 buffer[464] = 1;
 buffer[465] = 1;
 buffer[466] = 1;
 buffer[467] = 1;
 buffer[468] = 1;
 buffer[469] = 1;
 buffer[470] = 1;
 buffer[471] = 1;
 buffer[472] = 1;
 buffer[473] = 1;
 buffer[474] = 1;
 buffer[475] = 1;
 buffer[476] = 1;
 buffer[477] = 1;
 buffer[478] = 1;
 buffer[479] = 1;
 buffer[480] = 1;
 buffer[481] = 1;
 buffer[482] = 1;
 buffer[483] = 1;
 buffer[484] = 1;
 buffer[485] = 1;
 buffer[486] = 1;
 buffer[487] = 1;
 buffer[488] = 1;
 buffer[489] = 1;
 buffer[490] = 1;
 buffer[491] = 1;
 buffer[492] = 1;
 buffer[493] = 1;
 buffer[494] = 1;
 buffer[495] = 1;
 buffer[496] = 1;
 buffer[497] = 1;
 buffer[498] = 1;
 buffer[499] = 1;
 buffer[500] = 1;
 buffer[501] = 1;
 buffer[502] = 1;
 buffer[503] = 1;
 buffer[504] = 1;
 buffer[505] = 1;
 buffer[506] = 1;
 buffer[507] = 1;
 buffer[508] = 1;
 buffer[509] = 1;
 buffer[510] = 1;
 buffer[511] = 1;
end

endmodule

module M_apu_mem_waveformtable_2(
input                  [8:0] in_waveformtable_2_addr,
output reg  [3:0] out_waveformtable_2_rdata,
input                                   clock
);
reg  [3:0] buffer[511:0];
always @(posedge clock) begin
   out_waveformtable_2_rdata <= buffer[in_waveformtable_2_addr];
end
initial begin
 buffer[0] = 15;
 buffer[1] = 15;
 buffer[2] = 15;
 buffer[3] = 15;
 buffer[4] = 15;
 buffer[5] = 15;
 buffer[6] = 15;
 buffer[7] = 15;
 buffer[8] = 15;
 buffer[9] = 15;
 buffer[10] = 15;
 buffer[11] = 15;
 buffer[12] = 15;
 buffer[13] = 15;
 buffer[14] = 15;
 buffer[15] = 15;
 buffer[16] = 0;
 buffer[17] = 0;
 buffer[18] = 0;
 buffer[19] = 0;
 buffer[20] = 0;
 buffer[21] = 0;
 buffer[22] = 0;
 buffer[23] = 0;
 buffer[24] = 0;
 buffer[25] = 0;
 buffer[26] = 0;
 buffer[27] = 0;
 buffer[28] = 0;
 buffer[29] = 0;
 buffer[30] = 0;
 buffer[31] = 0;
 buffer[32] = 0;
 buffer[33] = 0;
 buffer[34] = 1;
 buffer[35] = 1;
 buffer[36] = 2;
 buffer[37] = 2;
 buffer[38] = 3;
 buffer[39] = 3;
 buffer[40] = 4;
 buffer[41] = 4;
 buffer[42] = 5;
 buffer[43] = 5;
 buffer[44] = 6;
 buffer[45] = 6;
 buffer[46] = 7;
 buffer[47] = 7;
 buffer[48] = 8;
 buffer[49] = 8;
 buffer[50] = 9;
 buffer[51] = 9;
 buffer[52] = 10;
 buffer[53] = 10;
 buffer[54] = 11;
 buffer[55] = 11;
 buffer[56] = 12;
 buffer[57] = 12;
 buffer[58] = 13;
 buffer[59] = 13;
 buffer[60] = 14;
 buffer[61] = 14;
 buffer[62] = 15;
 buffer[63] = 15;
 buffer[64] = 0;
 buffer[65] = 1;
 buffer[66] = 2;
 buffer[67] = 3;
 buffer[68] = 4;
 buffer[69] = 5;
 buffer[70] = 6;
 buffer[71] = 7;
 buffer[72] = 8;
 buffer[73] = 9;
 buffer[74] = 10;
 buffer[75] = 11;
 buffer[76] = 12;
 buffer[77] = 13;
 buffer[78] = 14;
 buffer[79] = 15;
 buffer[80] = 15;
 buffer[81] = 14;
 buffer[82] = 13;
 buffer[83] = 12;
 buffer[84] = 11;
 buffer[85] = 10;
 buffer[86] = 9;
 buffer[87] = 8;
 buffer[88] = 7;
 buffer[89] = 6;
 buffer[90] = 5;
 buffer[91] = 4;
 buffer[92] = 3;
 buffer[93] = 2;
 buffer[94] = 1;
 buffer[95] = 0;
 buffer[96] = 7;
 buffer[97] = 8;
 buffer[98] = 10;
 buffer[99] = 11;
 buffer[100] = 12;
 buffer[101] = 13;
 buffer[102] = 13;
 buffer[103] = 14;
 buffer[104] = 15;
 buffer[105] = 14;
 buffer[106] = 13;
 buffer[107] = 13;
 buffer[108] = 12;
 buffer[109] = 11;
 buffer[110] = 10;
 buffer[111] = 8;
 buffer[112] = 7;
 buffer[113] = 6;
 buffer[114] = 4;
 buffer[115] = 3;
 buffer[116] = 2;
 buffer[117] = 1;
 buffer[118] = 1;
 buffer[119] = 0;
 buffer[120] = 0;
 buffer[121] = 0;
 buffer[122] = 1;
 buffer[123] = 1;
 buffer[124] = 2;
 buffer[125] = 3;
 buffer[126] = 4;
 buffer[127] = 6;
 buffer[128] = 1;
 buffer[129] = 1;
 buffer[130] = 1;
 buffer[131] = 1;
 buffer[132] = 1;
 buffer[133] = 1;
 buffer[134] = 1;
 buffer[135] = 1;
 buffer[136] = 1;
 buffer[137] = 1;
 buffer[138] = 1;
 buffer[139] = 1;
 buffer[140] = 1;
 buffer[141] = 1;
 buffer[142] = 1;
 buffer[143] = 1;
 buffer[144] = 1;
 buffer[145] = 1;
 buffer[146] = 1;
 buffer[147] = 1;
 buffer[148] = 1;
 buffer[149] = 1;
 buffer[150] = 1;
 buffer[151] = 1;
 buffer[152] = 1;
 buffer[153] = 1;
 buffer[154] = 1;
 buffer[155] = 1;
 buffer[156] = 1;
 buffer[157] = 1;
 buffer[158] = 1;
 buffer[159] = 1;
 buffer[160] = 1;
 buffer[161] = 1;
 buffer[162] = 1;
 buffer[163] = 1;
 buffer[164] = 1;
 buffer[165] = 1;
 buffer[166] = 1;
 buffer[167] = 1;
 buffer[168] = 1;
 buffer[169] = 1;
 buffer[170] = 1;
 buffer[171] = 1;
 buffer[172] = 1;
 buffer[173] = 1;
 buffer[174] = 1;
 buffer[175] = 1;
 buffer[176] = 1;
 buffer[177] = 1;
 buffer[178] = 1;
 buffer[179] = 1;
 buffer[180] = 1;
 buffer[181] = 1;
 buffer[182] = 1;
 buffer[183] = 1;
 buffer[184] = 1;
 buffer[185] = 1;
 buffer[186] = 1;
 buffer[187] = 1;
 buffer[188] = 1;
 buffer[189] = 1;
 buffer[190] = 1;
 buffer[191] = 1;
 buffer[192] = 1;
 buffer[193] = 1;
 buffer[194] = 1;
 buffer[195] = 1;
 buffer[196] = 1;
 buffer[197] = 1;
 buffer[198] = 1;
 buffer[199] = 1;
 buffer[200] = 1;
 buffer[201] = 1;
 buffer[202] = 1;
 buffer[203] = 1;
 buffer[204] = 1;
 buffer[205] = 1;
 buffer[206] = 1;
 buffer[207] = 1;
 buffer[208] = 1;
 buffer[209] = 1;
 buffer[210] = 1;
 buffer[211] = 1;
 buffer[212] = 1;
 buffer[213] = 1;
 buffer[214] = 1;
 buffer[215] = 1;
 buffer[216] = 1;
 buffer[217] = 1;
 buffer[218] = 1;
 buffer[219] = 1;
 buffer[220] = 1;
 buffer[221] = 1;
 buffer[222] = 1;
 buffer[223] = 1;
 buffer[224] = 1;
 buffer[225] = 1;
 buffer[226] = 1;
 buffer[227] = 1;
 buffer[228] = 1;
 buffer[229] = 1;
 buffer[230] = 1;
 buffer[231] = 1;
 buffer[232] = 1;
 buffer[233] = 1;
 buffer[234] = 1;
 buffer[235] = 1;
 buffer[236] = 1;
 buffer[237] = 1;
 buffer[238] = 1;
 buffer[239] = 1;
 buffer[240] = 1;
 buffer[241] = 1;
 buffer[242] = 1;
 buffer[243] = 1;
 buffer[244] = 1;
 buffer[245] = 1;
 buffer[246] = 1;
 buffer[247] = 1;
 buffer[248] = 1;
 buffer[249] = 1;
 buffer[250] = 1;
 buffer[251] = 1;
 buffer[252] = 1;
 buffer[253] = 1;
 buffer[254] = 1;
 buffer[255] = 1;
 buffer[256] = 1;
 buffer[257] = 1;
 buffer[258] = 1;
 buffer[259] = 1;
 buffer[260] = 1;
 buffer[261] = 1;
 buffer[262] = 1;
 buffer[263] = 1;
 buffer[264] = 1;
 buffer[265] = 1;
 buffer[266] = 1;
 buffer[267] = 1;
 buffer[268] = 1;
 buffer[269] = 1;
 buffer[270] = 1;
 buffer[271] = 1;
 buffer[272] = 1;
 buffer[273] = 1;
 buffer[274] = 1;
 buffer[275] = 1;
 buffer[276] = 1;
 buffer[277] = 1;
 buffer[278] = 1;
 buffer[279] = 1;
 buffer[280] = 1;
 buffer[281] = 1;
 buffer[282] = 1;
 buffer[283] = 1;
 buffer[284] = 1;
 buffer[285] = 1;
 buffer[286] = 1;
 buffer[287] = 1;
 buffer[288] = 1;
 buffer[289] = 1;
 buffer[290] = 1;
 buffer[291] = 1;
 buffer[292] = 1;
 buffer[293] = 1;
 buffer[294] = 1;
 buffer[295] = 1;
 buffer[296] = 1;
 buffer[297] = 1;
 buffer[298] = 1;
 buffer[299] = 1;
 buffer[300] = 1;
 buffer[301] = 1;
 buffer[302] = 1;
 buffer[303] = 1;
 buffer[304] = 1;
 buffer[305] = 1;
 buffer[306] = 1;
 buffer[307] = 1;
 buffer[308] = 1;
 buffer[309] = 1;
 buffer[310] = 1;
 buffer[311] = 1;
 buffer[312] = 1;
 buffer[313] = 1;
 buffer[314] = 1;
 buffer[315] = 1;
 buffer[316] = 1;
 buffer[317] = 1;
 buffer[318] = 1;
 buffer[319] = 1;
 buffer[320] = 1;
 buffer[321] = 1;
 buffer[322] = 1;
 buffer[323] = 1;
 buffer[324] = 1;
 buffer[325] = 1;
 buffer[326] = 1;
 buffer[327] = 1;
 buffer[328] = 1;
 buffer[329] = 1;
 buffer[330] = 1;
 buffer[331] = 1;
 buffer[332] = 1;
 buffer[333] = 1;
 buffer[334] = 1;
 buffer[335] = 1;
 buffer[336] = 1;
 buffer[337] = 1;
 buffer[338] = 1;
 buffer[339] = 1;
 buffer[340] = 1;
 buffer[341] = 1;
 buffer[342] = 1;
 buffer[343] = 1;
 buffer[344] = 1;
 buffer[345] = 1;
 buffer[346] = 1;
 buffer[347] = 1;
 buffer[348] = 1;
 buffer[349] = 1;
 buffer[350] = 1;
 buffer[351] = 1;
 buffer[352] = 1;
 buffer[353] = 1;
 buffer[354] = 1;
 buffer[355] = 1;
 buffer[356] = 1;
 buffer[357] = 1;
 buffer[358] = 1;
 buffer[359] = 1;
 buffer[360] = 1;
 buffer[361] = 1;
 buffer[362] = 1;
 buffer[363] = 1;
 buffer[364] = 1;
 buffer[365] = 1;
 buffer[366] = 1;
 buffer[367] = 1;
 buffer[368] = 1;
 buffer[369] = 1;
 buffer[370] = 1;
 buffer[371] = 1;
 buffer[372] = 1;
 buffer[373] = 1;
 buffer[374] = 1;
 buffer[375] = 1;
 buffer[376] = 1;
 buffer[377] = 1;
 buffer[378] = 1;
 buffer[379] = 1;
 buffer[380] = 1;
 buffer[381] = 1;
 buffer[382] = 1;
 buffer[383] = 1;
 buffer[384] = 1;
 buffer[385] = 1;
 buffer[386] = 1;
 buffer[387] = 1;
 buffer[388] = 1;
 buffer[389] = 1;
 buffer[390] = 1;
 buffer[391] = 1;
 buffer[392] = 1;
 buffer[393] = 1;
 buffer[394] = 1;
 buffer[395] = 1;
 buffer[396] = 1;
 buffer[397] = 1;
 buffer[398] = 1;
 buffer[399] = 1;
 buffer[400] = 1;
 buffer[401] = 1;
 buffer[402] = 1;
 buffer[403] = 1;
 buffer[404] = 1;
 buffer[405] = 1;
 buffer[406] = 1;
 buffer[407] = 1;
 buffer[408] = 1;
 buffer[409] = 1;
 buffer[410] = 1;
 buffer[411] = 1;
 buffer[412] = 1;
 buffer[413] = 1;
 buffer[414] = 1;
 buffer[415] = 1;
 buffer[416] = 1;
 buffer[417] = 1;
 buffer[418] = 1;
 buffer[419] = 1;
 buffer[420] = 1;
 buffer[421] = 1;
 buffer[422] = 1;
 buffer[423] = 1;
 buffer[424] = 1;
 buffer[425] = 1;
 buffer[426] = 1;
 buffer[427] = 1;
 buffer[428] = 1;
 buffer[429] = 1;
 buffer[430] = 1;
 buffer[431] = 1;
 buffer[432] = 1;
 buffer[433] = 1;
 buffer[434] = 1;
 buffer[435] = 1;
 buffer[436] = 1;
 buffer[437] = 1;
 buffer[438] = 1;
 buffer[439] = 1;
 buffer[440] = 1;
 buffer[441] = 1;
 buffer[442] = 1;
 buffer[443] = 1;
 buffer[444] = 1;
 buffer[445] = 1;
 buffer[446] = 1;
 buffer[447] = 1;
 buffer[448] = 1;
 buffer[449] = 1;
 buffer[450] = 1;
 buffer[451] = 1;
 buffer[452] = 1;
 buffer[453] = 1;
 buffer[454] = 1;
 buffer[455] = 1;
 buffer[456] = 1;
 buffer[457] = 1;
 buffer[458] = 1;
 buffer[459] = 1;
 buffer[460] = 1;
 buffer[461] = 1;
 buffer[462] = 1;
 buffer[463] = 1;
 buffer[464] = 1;
 buffer[465] = 1;
 buffer[466] = 1;
 buffer[467] = 1;
 buffer[468] = 1;
 buffer[469] = 1;
 buffer[470] = 1;
 buffer[471] = 1;
 buffer[472] = 1;
 buffer[473] = 1;
 buffer[474] = 1;
 buffer[475] = 1;
 buffer[476] = 1;
 buffer[477] = 1;
 buffer[478] = 1;
 buffer[479] = 1;
 buffer[480] = 1;
 buffer[481] = 1;
 buffer[482] = 1;
 buffer[483] = 1;
 buffer[484] = 1;
 buffer[485] = 1;
 buffer[486] = 1;
 buffer[487] = 1;
 buffer[488] = 1;
 buffer[489] = 1;
 buffer[490] = 1;
 buffer[491] = 1;
 buffer[492] = 1;
 buffer[493] = 1;
 buffer[494] = 1;
 buffer[495] = 1;
 buffer[496] = 1;
 buffer[497] = 1;
 buffer[498] = 1;
 buffer[499] = 1;
 buffer[500] = 1;
 buffer[501] = 1;
 buffer[502] = 1;
 buffer[503] = 1;
 buffer[504] = 1;
 buffer[505] = 1;
 buffer[506] = 1;
 buffer[507] = 1;
 buffer[508] = 1;
 buffer[509] = 1;
 buffer[510] = 1;
 buffer[511] = 1;
end

endmodule

module M_apu_mem_frequencytable_1(
input                  [6:0] in_frequencytable_1_addr,
output reg  [15:0] out_frequencytable_1_rdata,
input                                   clock
);
reg  [15:0] buffer[127:0];
always @(posedge clock) begin
   out_frequencytable_1_rdata <= buffer[in_frequencytable_1_addr];
end
initial begin
 buffer[0] = 0;
 buffer[1] = 23889;
 buffer[2] = 22548;
 buffer[3] = 21283;
 buffer[4] = 20088;
 buffer[5] = 18961;
 buffer[6] = 17897;
 buffer[7] = 16892;
 buffer[8] = 15944;
 buffer[9] = 15049;
 buffer[10] = 14205;
 buffer[11] = 13407;
 buffer[12] = 12655;
 buffer[13] = 11945;
 buffer[14] = 11274;
 buffer[15] = 10641;
 buffer[16] = 10044;
 buffer[17] = 9480;
 buffer[18] = 8948;
 buffer[19] = 8446;
 buffer[20] = 7972;
 buffer[21] = 7525;
 buffer[22] = 7102;
 buffer[23] = 6704;
 buffer[24] = 6327;
 buffer[25] = 5972;
 buffer[26] = 5637;
 buffer[27] = 5321;
 buffer[28] = 5022;
 buffer[29] = 4740;
 buffer[30] = 4474;
 buffer[31] = 4223;
 buffer[32] = 3986;
 buffer[33] = 3762;
 buffer[34] = 3551;
 buffer[35] = 3352;
 buffer[36] = 3164;
 buffer[37] = 2896;
 buffer[38] = 2819;
 buffer[39] = 2660;
 buffer[40] = 2511;
 buffer[41] = 2370;
 buffer[42] = 2237;
 buffer[43] = 2112;
 buffer[44] = 1993;
 buffer[45] = 1881;
 buffer[46] = 1776;
 buffer[47] = 1676;
 buffer[48] = 1582;
 buffer[49] = 1493;
 buffer[50] = 1409;
 buffer[51] = 1330;
 buffer[52] = 1256;
 buffer[53] = 1185;
 buffer[54] = 1119;
 buffer[55] = 1056;
 buffer[56] = 997;
 buffer[57] = 941;
 buffer[58] = 888;
 buffer[59] = 838;
 buffer[60] = 791;
 buffer[61] = 747;
 buffer[62] = 705;
 buffer[63] = 665;
 buffer[64] = 1024;
 buffer[65] = 1024;
 buffer[66] = 1024;
 buffer[67] = 1024;
 buffer[68] = 1024;
 buffer[69] = 1024;
 buffer[70] = 1024;
 buffer[71] = 1024;
 buffer[72] = 1024;
 buffer[73] = 1024;
 buffer[74] = 1024;
 buffer[75] = 1024;
 buffer[76] = 1024;
 buffer[77] = 1024;
 buffer[78] = 1024;
 buffer[79] = 1024;
 buffer[80] = 1024;
 buffer[81] = 1024;
 buffer[82] = 1024;
 buffer[83] = 1024;
 buffer[84] = 1024;
 buffer[85] = 1024;
 buffer[86] = 1024;
 buffer[87] = 1024;
 buffer[88] = 1024;
 buffer[89] = 1024;
 buffer[90] = 1024;
 buffer[91] = 1024;
 buffer[92] = 1024;
 buffer[93] = 1024;
 buffer[94] = 1024;
 buffer[95] = 1024;
 buffer[96] = 1024;
 buffer[97] = 1024;
 buffer[98] = 1024;
 buffer[99] = 1024;
 buffer[100] = 1024;
 buffer[101] = 1024;
 buffer[102] = 1024;
 buffer[103] = 1024;
 buffer[104] = 1024;
 buffer[105] = 1024;
 buffer[106] = 1024;
 buffer[107] = 1024;
 buffer[108] = 1024;
 buffer[109] = 1024;
 buffer[110] = 1024;
 buffer[111] = 1024;
 buffer[112] = 1024;
 buffer[113] = 1024;
 buffer[114] = 1024;
 buffer[115] = 1024;
 buffer[116] = 1024;
 buffer[117] = 1024;
 buffer[118] = 1024;
 buffer[119] = 1024;
 buffer[120] = 1024;
 buffer[121] = 1024;
 buffer[122] = 1024;
 buffer[123] = 1024;
 buffer[124] = 1024;
 buffer[125] = 1024;
 buffer[126] = 1024;
 buffer[127] = 1024;
end

endmodule

module M_apu_mem_frequencytable_2(
input                  [6:0] in_frequencytable_2_addr,
output reg  [15:0] out_frequencytable_2_rdata,
input                                   clock
);
reg  [15:0] buffer[127:0];
always @(posedge clock) begin
   out_frequencytable_2_rdata <= buffer[in_frequencytable_2_addr];
end
initial begin
 buffer[0] = 0;
 buffer[1] = 23889;
 buffer[2] = 22548;
 buffer[3] = 21283;
 buffer[4] = 20088;
 buffer[5] = 18961;
 buffer[6] = 17897;
 buffer[7] = 16892;
 buffer[8] = 15944;
 buffer[9] = 15049;
 buffer[10] = 14205;
 buffer[11] = 13407;
 buffer[12] = 12655;
 buffer[13] = 11945;
 buffer[14] = 11274;
 buffer[15] = 10641;
 buffer[16] = 10044;
 buffer[17] = 9480;
 buffer[18] = 8948;
 buffer[19] = 8446;
 buffer[20] = 7972;
 buffer[21] = 7525;
 buffer[22] = 7102;
 buffer[23] = 6704;
 buffer[24] = 6327;
 buffer[25] = 5972;
 buffer[26] = 5637;
 buffer[27] = 5321;
 buffer[28] = 5022;
 buffer[29] = 4740;
 buffer[30] = 4474;
 buffer[31] = 4223;
 buffer[32] = 3986;
 buffer[33] = 3762;
 buffer[34] = 3551;
 buffer[35] = 3352;
 buffer[36] = 3164;
 buffer[37] = 2896;
 buffer[38] = 2819;
 buffer[39] = 2660;
 buffer[40] = 2511;
 buffer[41] = 2370;
 buffer[42] = 2237;
 buffer[43] = 2112;
 buffer[44] = 1993;
 buffer[45] = 1881;
 buffer[46] = 1776;
 buffer[47] = 1676;
 buffer[48] = 1582;
 buffer[49] = 1493;
 buffer[50] = 1409;
 buffer[51] = 1330;
 buffer[52] = 1256;
 buffer[53] = 1185;
 buffer[54] = 1119;
 buffer[55] = 1056;
 buffer[56] = 997;
 buffer[57] = 941;
 buffer[58] = 888;
 buffer[59] = 838;
 buffer[60] = 791;
 buffer[61] = 747;
 buffer[62] = 705;
 buffer[63] = 665;
 buffer[64] = 1024;
 buffer[65] = 1024;
 buffer[66] = 1024;
 buffer[67] = 1024;
 buffer[68] = 1024;
 buffer[69] = 1024;
 buffer[70] = 1024;
 buffer[71] = 1024;
 buffer[72] = 1024;
 buffer[73] = 1024;
 buffer[74] = 1024;
 buffer[75] = 1024;
 buffer[76] = 1024;
 buffer[77] = 1024;
 buffer[78] = 1024;
 buffer[79] = 1024;
 buffer[80] = 1024;
 buffer[81] = 1024;
 buffer[82] = 1024;
 buffer[83] = 1024;
 buffer[84] = 1024;
 buffer[85] = 1024;
 buffer[86] = 1024;
 buffer[87] = 1024;
 buffer[88] = 1024;
 buffer[89] = 1024;
 buffer[90] = 1024;
 buffer[91] = 1024;
 buffer[92] = 1024;
 buffer[93] = 1024;
 buffer[94] = 1024;
 buffer[95] = 1024;
 buffer[96] = 1024;
 buffer[97] = 1024;
 buffer[98] = 1024;
 buffer[99] = 1024;
 buffer[100] = 1024;
 buffer[101] = 1024;
 buffer[102] = 1024;
 buffer[103] = 1024;
 buffer[104] = 1024;
 buffer[105] = 1024;
 buffer[106] = 1024;
 buffer[107] = 1024;
 buffer[108] = 1024;
 buffer[109] = 1024;
 buffer[110] = 1024;
 buffer[111] = 1024;
 buffer[112] = 1024;
 buffer[113] = 1024;
 buffer[114] = 1024;
 buffer[115] = 1024;
 buffer[116] = 1024;
 buffer[117] = 1024;
 buffer[118] = 1024;
 buffer[119] = 1024;
 buffer[120] = 1024;
 buffer[121] = 1024;
 buffer[122] = 1024;
 buffer[123] = 1024;
 buffer[124] = 1024;
 buffer[125] = 1024;
 buffer[126] = 1024;
 buffer[127] = 1024;
end

endmodule

module M_apu (
in_waveform,
in_note,
in_duration,
in_apu_write,
in_staticGenerator,
out_audio_active,
out_audio_output,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [3:0] in_waveform;
input  [6:0] in_note;
input  [15:0] in_duration;
input  [1:0] in_apu_write;
input  [15:0] in_staticGenerator;
output  [0:0] out_audio_active;
output  [3:0] out_audio_output;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [3:0] _w_mem_waveformtable_1_rdata;
wire  [3:0] _w_mem_waveformtable_2_rdata;
wire  [15:0] _w_mem_frequencytable_1_rdata;
wire  [15:0] _w_mem_frequencytable_2_rdata;
reg  [15:0] _t_milliseconds_1;
reg  [15:0] _t_milliseconds_2;

reg  [8:0] _d_waveformtable_1_addr;
reg  [8:0] _q_waveformtable_1_addr;
reg  [8:0] _d_waveformtable_2_addr;
reg  [8:0] _q_waveformtable_2_addr;
reg  [6:0] _d_frequencytable_1_addr;
reg  [6:0] _q_frequencytable_1_addr;
reg  [6:0] _d_frequencytable_2_addr;
reg  [6:0] _q_frequencytable_2_addr;
reg  [2:0] _d_waveform_1;
reg  [2:0] _q_waveform_1;
reg  [5:0] _d_note_1;
reg  [5:0] _q_note_1;
reg  [4:0] _d_point_1;
reg  [4:0] _q_point_1;
reg  [15:0] _d_counter25mhz_1;
reg  [15:0] _q_counter25mhz_1;
reg  [15:0] _d_counter1khz_1;
reg  [15:0] _q_counter1khz_1;
reg  [2:0] _d_waveform_2;
reg  [2:0] _q_waveform_2;
reg  [5:0] _d_note_2;
reg  [5:0] _q_note_2;
reg  [4:0] _d_point_2;
reg  [4:0] _q_point_2;
reg  [15:0] _d_counter25mhz_2;
reg  [15:0] _q_counter25mhz_2;
reg  [15:0] _d_counter1khz_2;
reg  [15:0] _q_counter1khz_2;
reg  [15:0] _d_duration_1;
reg  [15:0] _q_duration_1;
reg  [15:0] _d_duration_2;
reg  [15:0] _q_duration_2;
reg  [0:0] _d_audio_active,_q_audio_active;
reg  [3:0] _d_audio_output,_q_audio_output;
reg  [1:0] _d_index,_q_index;
assign out_audio_active = _d_audio_active;
assign out_audio_output = _d_audio_output;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_waveformtable_1_addr <= 0;
_q_waveformtable_2_addr <= 0;
_q_frequencytable_1_addr <= 0;
_q_frequencytable_2_addr <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_waveformtable_1_addr <= _d_waveformtable_1_addr;
_q_waveformtable_2_addr <= _d_waveformtable_2_addr;
_q_frequencytable_1_addr <= _d_frequencytable_1_addr;
_q_frequencytable_2_addr <= _d_frequencytable_2_addr;
_q_waveform_1 <= _d_waveform_1;
_q_note_1 <= _d_note_1;
_q_point_1 <= _d_point_1;
_q_counter25mhz_1 <= _d_counter25mhz_1;
_q_counter1khz_1 <= _d_counter1khz_1;
_q_waveform_2 <= _d_waveform_2;
_q_note_2 <= _d_note_2;
_q_point_2 <= _d_point_2;
_q_counter25mhz_2 <= _d_counter25mhz_2;
_q_counter1khz_2 <= _d_counter1khz_2;
_q_duration_1 <= _d_duration_1;
_q_duration_2 <= _d_duration_2;
_q_audio_active <= _d_audio_active;
_q_audio_output <= _d_audio_output;
_q_index <= _d_index;
  end
end


M_apu_mem_waveformtable_1 __mem__waveformtable_1(
.clock(clock),
.in_waveformtable_1_addr(_d_waveformtable_1_addr),
.out_waveformtable_1_rdata(_w_mem_waveformtable_1_rdata)
);
M_apu_mem_waveformtable_2 __mem__waveformtable_2(
.clock(clock),
.in_waveformtable_2_addr(_d_waveformtable_2_addr),
.out_waveformtable_2_rdata(_w_mem_waveformtable_2_rdata)
);
M_apu_mem_frequencytable_1 __mem__frequencytable_1(
.clock(clock),
.in_frequencytable_1_addr(_d_frequencytable_1_addr),
.out_frequencytable_1_rdata(_w_mem_frequencytable_1_rdata)
);
M_apu_mem_frequencytable_2 __mem__frequencytable_2(
.clock(clock),
.in_frequencytable_2_addr(_d_frequencytable_2_addr),
.out_frequencytable_2_rdata(_w_mem_frequencytable_2_rdata)
);


always @* begin
_d_waveformtable_1_addr = _q_waveformtable_1_addr;
_d_waveformtable_2_addr = _q_waveformtable_2_addr;
_d_frequencytable_1_addr = _q_frequencytable_1_addr;
_d_frequencytable_2_addr = _q_frequencytable_2_addr;
_d_waveform_1 = _q_waveform_1;
_d_note_1 = _q_note_1;
_d_point_1 = _q_point_1;
_d_counter25mhz_1 = _q_counter25mhz_1;
_d_counter1khz_1 = _q_counter1khz_1;
_d_waveform_2 = _q_waveform_2;
_d_note_2 = _q_note_2;
_d_point_2 = _q_point_2;
_d_counter25mhz_2 = _q_counter25mhz_2;
_d_counter1khz_2 = _q_counter1khz_2;
_d_duration_1 = _q_duration_1;
_d_duration_2 = _q_duration_2;
_d_audio_active = _q_audio_active;
_d_audio_output = _q_audio_output;
_d_index = _q_index;
_t_milliseconds_1 = 0;
_t_milliseconds_2 = 0;
// _always_pre
_d_waveformtable_1_addr = _q_waveform_1*32+_q_point_1;
_d_waveformtable_2_addr = _q_waveform_2*32+_q_point_2;
_d_frequencytable_1_addr = _q_note_1;
_d_frequencytable_2_addr = _q_note_2;
_d_audio_active = (_q_duration_1>0)||(_q_duration_2>0);
if ((_q_duration_1!=0)&&(_q_counter25mhz_1==0)) begin
// __block_1
// __block_3
_d_audio_output = (_q_waveform_1==4)?in_staticGenerator:_w_mem_waveformtable_1_rdata;
// __block_4
end else begin
// __block_2
end
// __block_5
if ((_q_duration_2!=0)&&(_q_counter25mhz_2==0)) begin
// __block_6
// __block_8
_d_audio_output = (_q_waveform_2==4)?in_staticGenerator:_w_mem_waveformtable_2_rdata;
// __block_9
end else begin
// __block_7
end
// __block_10
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_waveformtable_1_addr = 0;
_d_waveformtable_2_addr = 0;
_d_frequencytable_1_addr = 0;
_d_frequencytable_2_addr = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_11
if (1) begin
// __block_12
// __block_14
  case (in_apu_write)
  1: begin
// __block_16_case
// __block_17
_d_waveform_1 = in_waveform;
_d_note_1 = in_note;
_d_duration_1 = in_duration;
_t_milliseconds_1 = 0;
_d_point_1 = 0;
_d_counter25mhz_1 = 0;
_d_counter1khz_1 = 25000;
// __block_18
  end
  2: begin
// __block_19_case
// __block_20
_d_waveform_2 = in_waveform;
_d_note_2 = in_note;
_d_duration_2 = in_duration;
_t_milliseconds_2 = 0;
_d_point_2 = 0;
_d_counter25mhz_2 = 0;
_d_counter1khz_2 = 25000;
// __block_21
  end
  default: begin
// __block_22_case
// __block_23
if (_q_duration_1!=0) begin
// __block_24
// __block_26
_d_counter25mhz_1 = (_q_counter25mhz_1!=0)?_q_counter25mhz_1-1:_w_mem_frequencytable_1_rdata;
_d_point_1 = (_d_counter25mhz_1!=0)?_q_point_1:_q_point_1+1;
_d_counter1khz_1 = (_q_counter1khz_1!=0)?_q_counter1khz_1-1:25000;
_d_duration_1 = (_d_counter1khz_1!=0)?_q_duration_1:_q_duration_1-1;
// __block_27
end else begin
// __block_25
end
// __block_28
if (_q_duration_2!=0) begin
// __block_29
// __block_31
_d_counter25mhz_2 = (_q_counter25mhz_2!=0)?_q_counter25mhz_2-1:_w_mem_frequencytable_2_rdata;
_d_point_2 = (_d_counter25mhz_2!=0)?_q_point_2:_q_point_2+1;
_d_counter1khz_2 = (_q_counter1khz_2!=0)?_q_counter1khz_2-1:25000;
_d_duration_2 = (_d_counter1khz_2!=0)?_q_duration_2:_q_duration_2-1;
// __block_32
end else begin
// __block_30
end
// __block_33
// __block_34
  end
endcase
// __block_15
// __block_35
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_13
_d_index = 3;
end
3: begin // end of apu
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_divmod32by16 (
in_dividendh,
in_dividendl,
in_divisor,
in_start,
out_quotient,
out_remainder,
out_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_dividendh;
input  [15:0] in_dividendl;
input  [15:0] in_divisor;
input  [1:0] in_start;
output  [15:0] out_quotient;
output  [15:0] out_remainder;
output  [0:0] out_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [31:0] _d_dividend_copy;
reg  [31:0] _q_dividend_copy;
reg  [31:0] _d_divisor_copy;
reg  [31:0] _q_divisor_copy;
reg  [31:0] _d_quotient_copy;
reg  [31:0] _q_quotient_copy;
reg  [31:0] _d_remainder_copy;
reg  [31:0] _q_remainder_copy;
reg  [0:0] _d_resultsign;
reg  [0:0] _q_resultsign;
reg  [5:0] _d_bit;
reg  [5:0] _q_bit;
reg  [15:0] _d_quotient,_q_quotient;
reg  [15:0] _d_remainder,_q_remainder;
reg  [0:0] _d_active,_q_active;
reg  [2:0] _d_index,_q_index;
assign out_quotient = _q_quotient;
assign out_remainder = _q_remainder;
assign out_active = _q_active;
assign out_done = (_q_index == 6);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_dividend_copy <= _d_dividend_copy;
_q_divisor_copy <= _d_divisor_copy;
_q_quotient_copy <= _d_quotient_copy;
_q_remainder_copy <= _d_remainder_copy;
_q_resultsign <= _d_resultsign;
_q_bit <= _d_bit;
_q_quotient <= _d_quotient;
_q_remainder <= _d_remainder;
_q_active <= _d_active;
_q_index <= _d_index;
  end
end




always @* begin
_d_dividend_copy = _q_dividend_copy;
_d_divisor_copy = _q_divisor_copy;
_d_quotient_copy = _q_quotient_copy;
_d_remainder_copy = _q_remainder_copy;
_d_resultsign = _q_resultsign;
_d_bit = _q_bit;
_d_quotient = _q_quotient;
_d_remainder = _q_remainder;
_d_active = _q_active;
_d_index = _q_index;
// _always_pre
_d_index = 6;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start!=0) begin
// __block_5
// __block_7
if (in_divisor==0) begin
// __block_8
// __block_10
_d_quotient_copy = 32'hffff;
_d_remainder_copy = in_divisor;
// __block_11
_d_index = 1;
end else begin
// __block_9
// __block_12
_d_bit = 32;
_d_quotient_copy = 0;
_d_remainder_copy = 0;
_d_dividend_copy = (in_start==1)?{in_dividendh,in_dividendl}:in_dividendh[15+:1]?-{in_dividendh,in_dividendl}:{in_dividendh,in_dividendl};
_d_divisor_copy = (in_start==1)?{16'b0,in_divisor}:in_divisor[15+:1]?{16'b0,-in_divisor}:{16'b0,in_divisor};
_d_resultsign = (in_start==1)?0:in_dividendh[15+:1]!=in_divisor[15+:1];
_d_active = 1;
_d_index = 3;
end
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_13
_d_index = 4;
end
2: begin
// __block_3
_d_index = 6;
end
4: begin
// __while__block_14
if (_q_bit!=0) begin
// __block_15
// __block_17
if ($unsigned({_q_remainder_copy[0+:31],_q_dividend_copy[_q_bit-1+:1]})>=$unsigned(_q_divisor_copy)) begin
// __block_18
// __block_20
_d_remainder_copy = {_q_remainder_copy[0+:31],_q_dividend_copy[_q_bit-1+:1]}-_q_divisor_copy;
_d_quotient_copy[_q_bit-1+:1] = 1;
// __block_21
end else begin
// __block_19
// __block_22
_d_remainder_copy = {_q_remainder_copy[0+:31],_q_dividend_copy[_q_bit-1+:1]};
// __block_23
end
// __block_24
_d_bit = _q_bit-1;
// __block_25
_d_index = 4;
end else begin
_d_index = 5;
end
end
5: begin
// __block_26
_d_quotient = _q_resultsign?-_q_quotient_copy[0+:16]:_q_quotient_copy[0+:16];
_d_remainder = _q_remainder_copy[0+:16];
_d_active = 0;
// __block_27
_d_index = 1;
end
6: begin // end of divmod32by16
end
default: begin 
_d_index = 6;
 end
endcase
end
endmodule


module M_divmod16by16 (
in_dividend,
in_divisor,
in_start,
out_quotient,
out_remainder,
out_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_dividend;
input  [15:0] in_divisor;
input  [0:0] in_start;
output  [15:0] out_quotient;
output  [15:0] out_remainder;
output  [0:0] out_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [15:0] _d_dividend_copy;
reg  [15:0] _q_dividend_copy;
reg  [15:0] _d_divisor_copy;
reg  [15:0] _q_divisor_copy;
reg  [15:0] _d_quotient_copy;
reg  [15:0] _q_quotient_copy;
reg  [15:0] _d_remainder_copy;
reg  [15:0] _q_remainder_copy;
reg  [0:0] _d_resultsign;
reg  [0:0] _q_resultsign;
reg  [5:0] _d_bit;
reg  [5:0] _q_bit;
reg  [15:0] _d_quotient,_q_quotient;
reg  [15:0] _d_remainder,_q_remainder;
reg  [0:0] _d_active,_q_active;
reg  [2:0] _d_index,_q_index;
assign out_quotient = _q_quotient;
assign out_remainder = _q_remainder;
assign out_active = _q_active;
assign out_done = (_q_index == 6);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_dividend_copy <= _d_dividend_copy;
_q_divisor_copy <= _d_divisor_copy;
_q_quotient_copy <= _d_quotient_copy;
_q_remainder_copy <= _d_remainder_copy;
_q_resultsign <= _d_resultsign;
_q_bit <= _d_bit;
_q_quotient <= _d_quotient;
_q_remainder <= _d_remainder;
_q_active <= _d_active;
_q_index <= _d_index;
  end
end




always @* begin
_d_dividend_copy = _q_dividend_copy;
_d_divisor_copy = _q_divisor_copy;
_d_quotient_copy = _q_quotient_copy;
_d_remainder_copy = _q_remainder_copy;
_d_resultsign = _q_resultsign;
_d_bit = _q_bit;
_d_quotient = _q_quotient;
_d_remainder = _q_remainder;
_d_active = _q_active;
_d_index = _q_index;
// _always_pre
_d_index = 6;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start) begin
// __block_5
// __block_7
if (in_divisor!=0) begin
// __block_8
// __block_10
_d_bit = 16;
_d_quotient_copy = 0;
_d_remainder_copy = 0;
_d_dividend_copy = in_dividend[15+:1]?-in_dividend:in_dividend;
_d_divisor_copy = in_divisor[15+:1]?-in_divisor:in_divisor;
_d_resultsign = in_dividend[15+:1]!=in_divisor[15+:1];
_d_active = 1;
_d_index = 3;
end else begin
// __block_9
// __block_26
_d_quotient_copy = 16'hffff;
_d_remainder_copy = in_divisor;
// __block_27
_d_index = 1;
end
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_11
_d_index = 4;
end
2: begin
// __block_3
_d_index = 6;
end
4: begin
// __while__block_12
if (_q_bit!=0) begin
// __block_13
// __block_15
if ($unsigned({_q_remainder_copy[0+:15],_q_dividend_copy[_q_bit-1+:1]})>=$unsigned(_q_divisor_copy)) begin
// __block_16
// __block_18
_d_remainder_copy = {_q_remainder_copy[0+:15],_q_dividend_copy[_q_bit-1+:1]}-_q_divisor_copy;
_d_quotient_copy[_q_bit-1+:1] = 1;
// __block_19
end else begin
// __block_17
// __block_20
_d_remainder_copy = {_q_remainder_copy[0+:15],_q_dividend_copy[_q_bit-1+:1]};
// __block_21
end
// __block_22
_d_bit = _q_bit-1;
// __block_23
_d_index = 4;
end else begin
_d_index = 5;
end
end
5: begin
// __block_24
_d_quotient = _q_resultsign?-_q_quotient_copy:_q_quotient_copy;
_d_remainder = _q_remainder_copy;
_d_active = 0;
// __block_25
_d_index = 1;
end
6: begin // end of divmod16by16
end
default: begin 
_d_index = 6;
 end
endcase
end
endmodule


module M_multi16by16to32DSP (
in_factor1,
in_factor2,
in_start,
out_product,
out_active,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_factor1;
input  [15:0] in_factor2;
input  [1:0] in_start;
output  [31:0] out_product;
output  [0:0] out_active;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [17:0] _d_factor1copy;
reg  [17:0] _q_factor1copy;
reg  [17:0] _d_factor2copy;
reg  [17:0] _q_factor2copy;
reg  [31:0] _d_nosignproduct;
reg  [31:0] _q_nosignproduct;
reg  [0:0] _d_productsign;
reg  [0:0] _q_productsign;
reg  [31:0] _d_product,_q_product;
reg  [0:0] _d_active,_q_active;
reg  [2:0] _d_index,_q_index;
assign out_product = _q_product;
assign out_active = _q_active;
assign out_done = (_q_index == 5);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_factor1copy <= _d_factor1copy;
_q_factor2copy <= _d_factor2copy;
_q_nosignproduct <= _d_nosignproduct;
_q_productsign <= _d_productsign;
_q_product <= _d_product;
_q_active <= _d_active;
_q_index <= _d_index;
  end
end




always @* begin
_d_factor1copy = _q_factor1copy;
_d_factor2copy = _q_factor2copy;
_d_nosignproduct = _q_nosignproduct;
_d_productsign = _q_productsign;
_d_product = _q_product;
_d_active = _q_active;
_d_index = _q_index;
// _always_pre
_d_index = 5;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (in_start!=0) begin
// __block_5
// __block_7
  case (in_start)
  1: begin
// __block_9_case
// __block_10
_d_factor1copy = in_factor1;
_d_factor2copy = in_factor2;
_d_productsign = 0;
// __block_11
  end
  2: begin
// __block_12_case
// __block_13
_d_product = 0;
_d_factor1copy = {2'b0,in_factor1[15+:1]?-in_factor1:in_factor1};
_d_factor2copy = {2'b0,in_factor2[15+:1]?-in_factor2:in_factor2};
_d_productsign = in_factor1[15+:1]!=in_factor2[15+:1];
// __block_14
  end
endcase
// __block_8
_d_product = 0;
_d_active = 1;
_d_index = 3;
end else begin
// __block_6
_d_index = 1;
end
end else begin
_d_index = 2;
end
end
3: begin
// __block_15
_d_nosignproduct = _q_factor1copy*_q_factor2copy;
_d_index = 4;
end
2: begin
// __block_3
_d_index = 5;
end
4: begin
// __block_16
_d_product = _q_productsign?-_q_nosignproduct:_q_nosignproduct;
_d_active = 0;
// __block_17
_d_index = 1;
end
5: begin // end of multi16by16to32DSP
end
default: begin 
_d_index = 5;
 end
endcase
end
endmodule


module M_doubleaddsub2input (
in_operand1h,
in_operand1l,
in_operand2h,
in_operand2l,
out_total,
out_difference,
out_binaryxor,
out_binaryor,
out_binaryand,
out_maximum,
out_minimum,
out_equal,
out_lessthan,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_operand1h;
input  [15:0] in_operand1l;
input  [15:0] in_operand2h;
input  [15:0] in_operand2l;
output  [31:0] out_total;
output  [31:0] out_difference;
output  [31:0] out_binaryxor;
output  [31:0] out_binaryor;
output  [31:0] out_binaryand;
output  [31:0] out_maximum;
output  [31:0] out_minimum;
output  [15:0] out_equal;
output  [15:0] out_lessthan;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [31:0] _w_operand1;
wire  [31:0] _w_operand2;

reg  [31:0] _d_total,_q_total;
reg  [31:0] _d_difference,_q_difference;
reg  [31:0] _d_binaryxor,_q_binaryxor;
reg  [31:0] _d_binaryor,_q_binaryor;
reg  [31:0] _d_binaryand,_q_binaryand;
reg  [31:0] _d_maximum,_q_maximum;
reg  [31:0] _d_minimum,_q_minimum;
reg  [15:0] _d_equal,_q_equal;
reg  [15:0] _d_lessthan,_q_lessthan;
reg  [1:0] _d_index,_q_index;
assign out_total = _q_total;
assign out_difference = _q_difference;
assign out_binaryxor = _q_binaryxor;
assign out_binaryor = _q_binaryor;
assign out_binaryand = _q_binaryand;
assign out_maximum = _q_maximum;
assign out_minimum = _q_minimum;
assign out_equal = _q_equal;
assign out_lessthan = _q_lessthan;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_total <= _d_total;
_q_difference <= _d_difference;
_q_binaryxor <= _d_binaryxor;
_q_binaryor <= _d_binaryor;
_q_binaryand <= _d_binaryand;
_q_maximum <= _d_maximum;
_q_minimum <= _d_minimum;
_q_equal <= _d_equal;
_q_lessthan <= _d_lessthan;
_q_index <= _d_index;
  end
end



assign _w_operand2 = {in_operand2h,in_operand2l};
assign _w_operand1 = {in_operand1h,in_operand1l};

always @* begin
_d_total = _q_total;
_d_difference = _q_difference;
_d_binaryxor = _q_binaryxor;
_d_binaryor = _q_binaryor;
_d_binaryand = _q_binaryand;
_d_maximum = _q_maximum;
_d_minimum = _q_minimum;
_d_equal = _q_equal;
_d_lessthan = _q_lessthan;
_d_index = _q_index;
// _always_pre
_d_total = _w_operand1+_w_operand2;
_d_difference = _w_operand1-_w_operand2;
_d_binaryxor = _w_operand1^_w_operand2;
_d_binaryor = _w_operand1|_w_operand2;
_d_binaryand = _w_operand1&_w_operand2;
_d_maximum = (_w_operand1>_w_operand2)?_w_operand1:_w_operand2;
_d_minimum = (_w_operand1<_w_operand2)?_w_operand1:_w_operand2;
_d_equal = {16{(_w_operand1==_w_operand2)}};
_d_lessthan = {16{(_w_operand1<_w_operand2)}};
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
// __block_5
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of doubleaddsub2input
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_doubleaddsub1input (
in_operand1h,
in_operand1l,
out_increment,
out_decrement,
out_times2,
out_divide2,
out_negation,
out_binaryinvert,
out_absolute,
out_zeroequal,
out_zeroless,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_operand1h;
input  [15:0] in_operand1l;
output  [31:0] out_increment;
output  [31:0] out_decrement;
output  [31:0] out_times2;
output  [31:0] out_divide2;
output  [31:0] out_negation;
output  [31:0] out_binaryinvert;
output  [31:0] out_absolute;
output  [15:0] out_zeroequal;
output  [15:0] out_zeroless;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [31:0] _w_operand1;

reg  [31:0] _d_increment,_q_increment;
reg  [31:0] _d_decrement,_q_decrement;
reg  [31:0] _d_times2,_q_times2;
reg  [31:0] _d_divide2,_q_divide2;
reg  [31:0] _d_negation,_q_negation;
reg  [31:0] _d_binaryinvert,_q_binaryinvert;
reg  [31:0] _d_absolute,_q_absolute;
reg  [15:0] _d_zeroequal,_q_zeroequal;
reg  [15:0] _d_zeroless,_q_zeroless;
reg  [1:0] _d_index,_q_index;
assign out_increment = _q_increment;
assign out_decrement = _q_decrement;
assign out_times2 = _q_times2;
assign out_divide2 = _q_divide2;
assign out_negation = _q_negation;
assign out_binaryinvert = _q_binaryinvert;
assign out_absolute = _q_absolute;
assign out_zeroequal = _q_zeroequal;
assign out_zeroless = _q_zeroless;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_increment <= _d_increment;
_q_decrement <= _d_decrement;
_q_times2 <= _d_times2;
_q_divide2 <= _d_divide2;
_q_negation <= _d_negation;
_q_binaryinvert <= _d_binaryinvert;
_q_absolute <= _d_absolute;
_q_zeroequal <= _d_zeroequal;
_q_zeroless <= _d_zeroless;
_q_index <= _d_index;
  end
end



assign _w_operand1 = {in_operand1h,in_operand1l};

always @* begin
_d_increment = _q_increment;
_d_decrement = _q_decrement;
_d_times2 = _q_times2;
_d_divide2 = _q_divide2;
_d_negation = _q_negation;
_d_binaryinvert = _q_binaryinvert;
_d_absolute = _q_absolute;
_d_zeroequal = _q_zeroequal;
_d_zeroless = _q_zeroless;
_d_index = _q_index;
// _always_pre
_d_increment = _w_operand1+1;
_d_decrement = _w_operand1-1;
_d_times2 = _w_operand1<<1;
_d_divide2 = {_w_operand1[31+:1],_w_operand1[1+:31]};
_d_negation = -_w_operand1;
_d_binaryinvert = ~_w_operand1;
_d_absolute = (_w_operand1[31+:1])?-_w_operand1:_w_operand1;
_d_zeroequal = {16{(_w_operand1==0)}};
_d_zeroless = {16{(_w_operand1<0)}};
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
// __block_5
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of doubleaddsub1input
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_memmap_io_mem_bitmap(
input      [18:0]                in_bitmap_addr0,
output reg  [6:0]     out_bitmap_rdata0,
output reg  [6:0]     out_bitmap_rdata1,
input      [0:0]             in_bitmap_wenable1,
input      [6:0]                 in_bitmap_wdata1,
input      [18:0]                in_bitmap_addr1,
input      clock0,
input      clock1
);
reg  [6:0] buffer[307199:0];
always @(posedge clock0) begin
  out_bitmap_rdata0 <= buffer[in_bitmap_addr0];
end
always @(posedge clock1) begin
  if (in_bitmap_wenable1) begin
    buffer[in_bitmap_addr1] <= in_bitmap_wdata1;
  end
end

endmodule

module M_memmap_io_mem_uartInBuffer(
input      [11:0]                in_uartInBuffer_addr0,
output reg  [7:0]     out_uartInBuffer_rdata0,
output reg  [7:0]     out_uartInBuffer_rdata1,
input      [0:0]             in_uartInBuffer_wenable1,
input      [7:0]                 in_uartInBuffer_wdata1,
input      [11:0]                in_uartInBuffer_addr1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[4095:0];
always @(posedge clock0) begin
  out_uartInBuffer_rdata0 <= buffer[in_uartInBuffer_addr0];
end
always @(posedge clock1) begin
  if (in_uartInBuffer_wenable1) begin
    buffer[in_uartInBuffer_addr1] <= in_uartInBuffer_wdata1;
  end
end

endmodule

module M_memmap_io_mem_uartOutBuffer(
input      [7:0]                in_uartOutBuffer_addr0,
output reg  [7:0]     out_uartOutBuffer_rdata0,
output reg  [7:0]     out_uartOutBuffer_rdata1,
input      [0:0]             in_uartOutBuffer_wenable1,
input      [7:0]                 in_uartOutBuffer_wdata1,
input      [7:0]                in_uartOutBuffer_addr1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[255:0];
always @(posedge clock0) begin
  out_uartOutBuffer_rdata0 <= buffer[in_uartOutBuffer_addr0];
end
always @(posedge clock1) begin
  if (in_uartOutBuffer_wenable1) begin
    buffer[in_uartOutBuffer_addr1] <= in_uartOutBuffer_wdata1;
  end
end

endmodule

module M_memmap_io (
in_btns,
in_uart_rx,
in_vblank,
in_pix_active,
in_pix_x,
in_pix_y,
in_clock_50mhz,
in_clock_25mhz,
in_video_clock,
in_video_reset,
in_memoryAddress,
in_writeData,
in_memoryWrite,
in_memoryRead,
out_leds,
out_uart_tx,
out_audio_l,
out_audio_r,
out_video_r,
out_video_g,
out_video_b,
out_readData,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [6:0] in_btns;
input  [0:0] in_uart_rx;
input  [0:0] in_vblank;
input  [0:0] in_pix_active;
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_clock_50mhz;
input  [0:0] in_clock_25mhz;
input  [0:0] in_video_clock;
input  [0:0] in_video_reset;
input  [15:0] in_memoryAddress;
input  [15:0] in_writeData;
input  [0:0] in_memoryWrite;
input  [0:0] in_memoryRead;
output  [7:0] out_leds;
output  [0:0] out_uart_tx;
output  [3:0] out_audio_l;
output  [3:0] out_audio_r;
output  [7:0] out_video_r;
output  [7:0] out_video_g;
output  [7:0] out_video_b;
output  [15:0] out_readData;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [15:0] _w_p1hz_counter1hz;
wire _w_p1hz_done;
wire  [15:0] _w_timer1hz_counter1hz;
wire _w_timer1hz_done;
wire  [15:0] _w_sleepTimer_counter1khz;
wire _w_sleepTimer_done;
wire  [15:0] _w_timer1khz_counter1khz;
wire _w_timer1khz_done;
wire  [15:0] _w_rng_g_noise_out;
wire  [15:0] _w_rng_u_noise_out;
wire _w_rng_done;
wire  [0:0] _w_usend_io_busy;
wire  [0:0] _w_usend_uart_tx;
wire _w_usend_done;
wire  [7:0] _w_urecv_io_data_out;
wire  [0:0] _w_urecv_io_data_out_ready;
wire  [1:0] _w_background_generator_pix_red;
wire  [1:0] _w_background_generator_pix_green;
wire  [1:0] _w_background_generator_pix_blue;
wire _w_background_generator_done;
wire  [1:0] _w_tile_map_pix_red;
wire  [1:0] _w_tile_map_pix_green;
wire  [1:0] _w_tile_map_pix_blue;
wire  [0:0] _w_tile_map_tilemap_display;
wire  [3:0] _w_tile_map_tm_lastaction;
wire  [1:0] _w_tile_map_tm_active;
wire _w_tile_map_done;
wire  [1:0] _w_bitmap_window_pix_red;
wire  [1:0] _w_bitmap_window_pix_green;
wire  [1:0] _w_bitmap_window_pix_blue;
wire  [0:0] _w_bitmap_window_bitmap_display;
wire  [9:0] _w_bitmap_window_x_offset;
wire  [9:0] _w_bitmap_window_y_offset;
wire  [6:0] _w_bitmap_window_bitmap_colour_read;
wire  [18:0] _w_bitmap_window_bitmap_addr0;
wire _w_bitmap_window_done;
wire  [18:0] _w_pixel_writer_bitmap_addr1;
wire  [0:0] _w_pixel_writer_bitmap_wenable1;
wire  [6:0] _w_pixel_writer_bitmap_wdata1;
wire _w_pixel_writer_done;
wire  [1:0] _w_lower_sprites_pix_red;
wire  [1:0] _w_lower_sprites_pix_green;
wire  [1:0] _w_lower_sprites_pix_blue;
wire  [0:0] _w_lower_sprites_sprite_layer_display;
wire  [0:0] _w_lower_sprites_sprite_read_active;
wire  [0:0] _w_lower_sprites_sprite_read_double;
wire  [5:0] _w_lower_sprites_sprite_read_colour;
wire signed [10:0] _w_lower_sprites_sprite_read_x;
wire signed [10:0] _w_lower_sprites_sprite_read_y;
wire  [2:0] _w_lower_sprites_sprite_read_tile;
wire  [15:0] _w_lower_sprites_collision_0;
wire  [15:0] _w_lower_sprites_collision_1;
wire  [15:0] _w_lower_sprites_collision_2;
wire  [15:0] _w_lower_sprites_collision_3;
wire  [15:0] _w_lower_sprites_collision_4;
wire  [15:0] _w_lower_sprites_collision_5;
wire  [15:0] _w_lower_sprites_collision_6;
wire  [15:0] _w_lower_sprites_collision_7;
wire  [15:0] _w_lower_sprites_collision_8;
wire  [15:0] _w_lower_sprites_collision_9;
wire  [15:0] _w_lower_sprites_collision_10;
wire  [15:0] _w_lower_sprites_collision_11;
wire  [15:0] _w_lower_sprites_collision_12;
wire _w_lower_sprites_done;
wire  [1:0] _w_upper_sprites_pix_red;
wire  [1:0] _w_upper_sprites_pix_green;
wire  [1:0] _w_upper_sprites_pix_blue;
wire  [0:0] _w_upper_sprites_sprite_layer_display;
wire  [0:0] _w_upper_sprites_sprite_read_active;
wire  [0:0] _w_upper_sprites_sprite_read_double;
wire  [5:0] _w_upper_sprites_sprite_read_colour;
wire signed [10:0] _w_upper_sprites_sprite_read_x;
wire signed [10:0] _w_upper_sprites_sprite_read_y;
wire  [2:0] _w_upper_sprites_sprite_read_tile;
wire  [15:0] _w_upper_sprites_collision_0;
wire  [15:0] _w_upper_sprites_collision_1;
wire  [15:0] _w_upper_sprites_collision_2;
wire  [15:0] _w_upper_sprites_collision_3;
wire  [15:0] _w_upper_sprites_collision_4;
wire  [15:0] _w_upper_sprites_collision_5;
wire  [15:0] _w_upper_sprites_collision_6;
wire  [15:0] _w_upper_sprites_collision_7;
wire  [15:0] _w_upper_sprites_collision_8;
wire  [15:0] _w_upper_sprites_collision_9;
wire  [15:0] _w_upper_sprites_collision_10;
wire  [15:0] _w_upper_sprites_collision_11;
wire  [15:0] _w_upper_sprites_collision_12;
wire _w_upper_sprites_done;
wire  [1:0] _w_character_map_window_pix_red;
wire  [1:0] _w_character_map_window_pix_green;
wire  [1:0] _w_character_map_window_pix_blue;
wire  [0:0] _w_character_map_window_character_map_display;
wire  [0:0] _w_character_map_window_tpu_active;
wire _w_character_map_window_done;
wire  [1:0] _w_terminal_window_pix_red;
wire  [1:0] _w_terminal_window_pix_green;
wire  [1:0] _w_terminal_window_pix_blue;
wire  [0:0] _w_terminal_window_terminal_display;
wire  [1:0] _w_terminal_window_terminal_active;
wire _w_terminal_window_done;
wire  [7:0] _w_display_pix_red;
wire  [7:0] _w_display_pix_green;
wire  [7:0] _w_display_pix_blue;
wire _w_display_done;
wire  [0:0] _w_apu_processor_L_audio_active;
wire  [3:0] _w_apu_processor_L_audio_output;
wire _w_apu_processor_L_done;
wire  [0:0] _w_apu_processor_R_audio_active;
wire  [3:0] _w_apu_processor_R_audio_output;
wire _w_apu_processor_R_done;
wire signed [10:0] _w_gpu_processor_bitmap_x_write;
wire signed [10:0] _w_gpu_processor_bitmap_y_write;
wire  [6:0] _w_gpu_processor_bitmap_colour_write;
wire  [0:0] _w_gpu_processor_bitmap_write;
wire  [0:0] _w_gpu_processor_gpu_active;
wire  [0:0] _w_gpu_processor_vector_block_active;
wire _w_gpu_processor_done;
wire  [15:0] _w_divmod32by16to16qr_quotient;
wire  [15:0] _w_divmod32by16to16qr_remainder;
wire  [0:0] _w_divmod32by16to16qr_active;
wire _w_divmod32by16to16qr_done;
wire  [15:0] _w_divmod16by16to16qr_quotient;
wire  [15:0] _w_divmod16by16to16qr_remainder;
wire  [0:0] _w_divmod16by16to16qr_active;
wire _w_divmod16by16to16qr_done;
wire  [31:0] _w_multiplier16by16to32_product;
wire  [0:0] _w_multiplier16by16to32_active;
wire _w_multiplier16by16to32_done;
wire  [31:0] _w_doperations2_total;
wire  [31:0] _w_doperations2_difference;
wire  [31:0] _w_doperations2_binaryxor;
wire  [31:0] _w_doperations2_binaryor;
wire  [31:0] _w_doperations2_binaryand;
wire  [31:0] _w_doperations2_maximum;
wire  [31:0] _w_doperations2_minimum;
wire  [15:0] _w_doperations2_equal;
wire  [15:0] _w_doperations2_lessthan;
wire _w_doperations2_done;
wire  [31:0] _w_doperations1_increment;
wire  [31:0] _w_doperations1_decrement;
wire  [31:0] _w_doperations1_times2;
wire  [31:0] _w_doperations1_divide2;
wire  [31:0] _w_doperations1_negation;
wire  [31:0] _w_doperations1_binaryinvert;
wire  [31:0] _w_doperations1_absolute;
wire  [15:0] _w_doperations1_zeroequal;
wire  [15:0] _w_doperations1_zeroless;
wire _w_doperations1_done;
wire  [6:0] _w_mem_bitmap_rdata0;
wire  [7:0] _w_mem_uartInBuffer_rdata0;
wire  [7:0] _w_mem_uartOutBuffer_rdata0;
reg  [6:0] _t_reg_btns;

reg  [7:0] _d_uo_data_in;
reg  [7:0] _q_uo_data_in;
reg  [0:0] _d_uo_data_in_ready;
reg  [0:0] _q_uo_data_in_ready;
reg  [11:0] _d_uartInBuffer_addr0;
reg  [11:0] _q_uartInBuffer_addr0;
reg  [0:0] _d_uartInBuffer_wenable1;
reg  [0:0] _q_uartInBuffer_wenable1;
reg  [7:0] _d_uartInBuffer_wdata1;
reg  [7:0] _q_uartInBuffer_wdata1;
reg  [11:0] _d_uartInBuffer_addr1;
reg  [11:0] _q_uartInBuffer_addr1;
reg  [12:0] _d_uartInBufferNext;
reg  [12:0] _q_uartInBufferNext;
reg  [12:0] _d_uartInBufferTop;
reg  [12:0] _q_uartInBufferTop;
reg  [7:0] _d_uartOutBuffer_addr0;
reg  [7:0] _q_uartOutBuffer_addr0;
reg  [0:0] _d_uartOutBuffer_wenable1;
reg  [0:0] _q_uartOutBuffer_wenable1;
reg  [7:0] _d_uartOutBuffer_wdata1;
reg  [7:0] _q_uartOutBuffer_wdata1;
reg  [7:0] _d_uartOutBuffer_addr1;
reg  [7:0] _q_uartOutBuffer_addr1;
reg  [7:0] _d_uartOutBufferNext;
reg  [7:0] _q_uartOutBufferNext;
reg  [7:0] _d_uartOutBufferTop;
reg  [7:0] _q_uartOutBufferTop;
reg  [7:0] _d_newuartOutBufferTop;
reg  [7:0] _q_newuartOutBufferTop;
reg  [1:0] _d_coProReset;
reg  [1:0] _q_coProReset;
reg  [6:0] _d_delayed_4582_4;
reg  [6:0] _q_delayed_4582_4;
reg  [7:0] _d_leds,_q_leds;
reg  [15:0] _d_readData,_q_readData;
reg  [0:0] _d_p1hz_resetCounter,_q_p1hz_resetCounter;
reg  [0:0] _d_timer1hz_resetCounter,_q_timer1hz_resetCounter;
reg  [15:0] _d_sleepTimer_resetCount,_q_sleepTimer_resetCount;
reg  [0:0] _d_sleepTimer_resetCounter,_q_sleepTimer_resetCounter;
reg  [15:0] _d_timer1khz_resetCount,_q_timer1khz_resetCount;
reg  [0:0] _d_timer1khz_resetCounter,_q_timer1khz_resetCounter;
reg  [0:0] _d_rng_resetRandom,_q_rng_resetRandom;
reg  [5:0] _d_background_generator_backgroundcolour,_q_background_generator_backgroundcolour;
reg  [5:0] _d_background_generator_backgroundcolour_alt,_q_background_generator_backgroundcolour_alt;
reg  [3:0] _d_background_generator_backgroundcolour_mode,_q_background_generator_backgroundcolour_mode;
reg  [2:0] _d_background_generator_background_write,_q_background_generator_background_write;
reg  [5:0] _d_tile_map_tm_x,_q_tile_map_tm_x;
reg  [5:0] _d_tile_map_tm_y,_q_tile_map_tm_y;
reg  [4:0] _d_tile_map_tm_character,_q_tile_map_tm_character;
reg  [5:0] _d_tile_map_tm_foreground,_q_tile_map_tm_foreground;
reg  [6:0] _d_tile_map_tm_background,_q_tile_map_tm_background;
reg  [0:0] _d_tile_map_tm_write,_q_tile_map_tm_write;
reg  [4:0] _d_tile_map_tile_writer_tile,_q_tile_map_tile_writer_tile;
reg  [3:0] _d_tile_map_tile_writer_line,_q_tile_map_tile_writer_line;
reg  [15:0] _d_tile_map_tile_writer_bitmap,_q_tile_map_tile_writer_bitmap;
reg  [3:0] _d_tile_map_tm_scrollwrap,_q_tile_map_tm_scrollwrap;
reg  [2:0] _d_bitmap_window_bitmap_write_offset,_q_bitmap_window_bitmap_write_offset;
reg signed [15:0] _d_bitmap_window_bitmap_x_read,_q_bitmap_window_bitmap_x_read;
reg signed [15:0] _d_bitmap_window_bitmap_y_read,_q_bitmap_window_bitmap_y_read;
reg  [3:0] _d_lower_sprites_sprite_set_number,_q_lower_sprites_sprite_set_number;
reg  [0:0] _d_lower_sprites_sprite_set_active,_q_lower_sprites_sprite_set_active;
reg  [0:0] _d_lower_sprites_sprite_set_double,_q_lower_sprites_sprite_set_double;
reg  [5:0] _d_lower_sprites_sprite_set_colour,_q_lower_sprites_sprite_set_colour;
reg signed [10:0] _d_lower_sprites_sprite_set_x,_q_lower_sprites_sprite_set_x;
reg signed [10:0] _d_lower_sprites_sprite_set_y,_q_lower_sprites_sprite_set_y;
reg  [2:0] _d_lower_sprites_sprite_set_tile,_q_lower_sprites_sprite_set_tile;
reg  [3:0] _d_lower_sprites_sprite_layer_write,_q_lower_sprites_sprite_layer_write;
reg  [15:0] _d_lower_sprites_sprite_update,_q_lower_sprites_sprite_update;
reg  [3:0] _d_lower_sprites_sprite_writer_sprite,_q_lower_sprites_sprite_writer_sprite;
reg  [6:0] _d_lower_sprites_sprite_writer_line,_q_lower_sprites_sprite_writer_line;
reg  [15:0] _d_lower_sprites_sprite_writer_bitmap,_q_lower_sprites_sprite_writer_bitmap;
reg  [0:0] _d_lower_sprites_sprite_writer_active,_q_lower_sprites_sprite_writer_active;
reg  [3:0] _d_upper_sprites_sprite_set_number,_q_upper_sprites_sprite_set_number;
reg  [0:0] _d_upper_sprites_sprite_set_active,_q_upper_sprites_sprite_set_active;
reg  [0:0] _d_upper_sprites_sprite_set_double,_q_upper_sprites_sprite_set_double;
reg  [5:0] _d_upper_sprites_sprite_set_colour,_q_upper_sprites_sprite_set_colour;
reg signed [10:0] _d_upper_sprites_sprite_set_x,_q_upper_sprites_sprite_set_x;
reg signed [10:0] _d_upper_sprites_sprite_set_y,_q_upper_sprites_sprite_set_y;
reg  [2:0] _d_upper_sprites_sprite_set_tile,_q_upper_sprites_sprite_set_tile;
reg  [3:0] _d_upper_sprites_sprite_layer_write,_q_upper_sprites_sprite_layer_write;
reg  [15:0] _d_upper_sprites_sprite_update,_q_upper_sprites_sprite_update;
reg  [3:0] _d_upper_sprites_sprite_writer_sprite,_q_upper_sprites_sprite_writer_sprite;
reg  [6:0] _d_upper_sprites_sprite_writer_line,_q_upper_sprites_sprite_writer_line;
reg  [15:0] _d_upper_sprites_sprite_writer_bitmap,_q_upper_sprites_sprite_writer_bitmap;
reg  [0:0] _d_upper_sprites_sprite_writer_active,_q_upper_sprites_sprite_writer_active;
reg  [6:0] _d_character_map_window_tpu_x,_q_character_map_window_tpu_x;
reg  [4:0] _d_character_map_window_tpu_y,_q_character_map_window_tpu_y;
reg  [7:0] _d_character_map_window_tpu_character,_q_character_map_window_tpu_character;
reg  [5:0] _d_character_map_window_tpu_foreground,_q_character_map_window_tpu_foreground;
reg  [6:0] _d_character_map_window_tpu_background,_q_character_map_window_tpu_background;
reg  [2:0] _d_character_map_window_tpu_write,_q_character_map_window_tpu_write;
reg  [7:0] _d_terminal_window_terminal_character,_q_terminal_window_terminal_character;
reg  [1:0] _d_terminal_window_terminal_write,_q_terminal_window_terminal_write;
reg  [0:0] _d_terminal_window_showterminal,_q_terminal_window_showterminal;
reg  [3:0] _d_apu_processor_L_waveform,_q_apu_processor_L_waveform;
reg  [6:0] _d_apu_processor_L_note,_q_apu_processor_L_note;
reg  [15:0] _d_apu_processor_L_duration,_q_apu_processor_L_duration;
reg  [1:0] _d_apu_processor_L_apu_write,_q_apu_processor_L_apu_write;
reg  [3:0] _d_apu_processor_R_waveform,_q_apu_processor_R_waveform;
reg  [6:0] _d_apu_processor_R_note,_q_apu_processor_R_note;
reg  [15:0] _d_apu_processor_R_duration,_q_apu_processor_R_duration;
reg  [1:0] _d_apu_processor_R_apu_write,_q_apu_processor_R_apu_write;
reg signed [10:0] _d_gpu_processor_gpu_x,_q_gpu_processor_gpu_x;
reg signed [10:0] _d_gpu_processor_gpu_y,_q_gpu_processor_gpu_y;
reg  [7:0] _d_gpu_processor_gpu_colour,_q_gpu_processor_gpu_colour;
reg signed [10:0] _d_gpu_processor_gpu_param0,_q_gpu_processor_gpu_param0;
reg signed [10:0] _d_gpu_processor_gpu_param1,_q_gpu_processor_gpu_param1;
reg signed [10:0] _d_gpu_processor_gpu_param2,_q_gpu_processor_gpu_param2;
reg signed [10:0] _d_gpu_processor_gpu_param3,_q_gpu_processor_gpu_param3;
reg  [3:0] _d_gpu_processor_gpu_write,_q_gpu_processor_gpu_write;
reg  [4:0] _d_gpu_processor_blit1_writer_tile,_q_gpu_processor_blit1_writer_tile;
reg  [3:0] _d_gpu_processor_blit1_writer_line,_q_gpu_processor_blit1_writer_line;
reg  [15:0] _d_gpu_processor_blit1_writer_bitmap,_q_gpu_processor_blit1_writer_bitmap;
reg  [4:0] _d_gpu_processor_vector_block_number,_q_gpu_processor_vector_block_number;
reg  [6:0] _d_gpu_processor_vector_block_colour,_q_gpu_processor_vector_block_colour;
reg signed [10:0] _d_gpu_processor_vector_block_xc,_q_gpu_processor_vector_block_xc;
reg signed [10:0] _d_gpu_processor_vector_block_yc,_q_gpu_processor_vector_block_yc;
reg  [0:0] _d_gpu_processor_draw_vector,_q_gpu_processor_draw_vector;
reg  [4:0] _d_gpu_processor_vertices_writer_block,_q_gpu_processor_vertices_writer_block;
reg  [5:0] _d_gpu_processor_vertices_writer_vertex,_q_gpu_processor_vertices_writer_vertex;
reg signed [5:0] _d_gpu_processor_vertices_writer_xdelta,_q_gpu_processor_vertices_writer_xdelta;
reg signed [5:0] _d_gpu_processor_vertices_writer_ydelta,_q_gpu_processor_vertices_writer_ydelta;
reg  [0:0] _d_gpu_processor_vertices_writer_active,_q_gpu_processor_vertices_writer_active;
reg  [15:0] _d_divmod32by16to16qr_dividendh,_q_divmod32by16to16qr_dividendh;
reg  [15:0] _d_divmod32by16to16qr_dividendl,_q_divmod32by16to16qr_dividendl;
reg  [15:0] _d_divmod32by16to16qr_divisor,_q_divmod32by16to16qr_divisor;
reg  [1:0] _d_divmod32by16to16qr_start,_q_divmod32by16to16qr_start;
reg  [15:0] _d_divmod16by16to16qr_dividend,_q_divmod16by16to16qr_dividend;
reg  [15:0] _d_divmod16by16to16qr_divisor,_q_divmod16by16to16qr_divisor;
reg  [0:0] _d_divmod16by16to16qr_start,_q_divmod16by16to16qr_start;
reg  [15:0] _d_multiplier16by16to32_factor1,_q_multiplier16by16to32_factor1;
reg  [15:0] _d_multiplier16by16to32_factor2,_q_multiplier16by16to32_factor2;
reg  [1:0] _d_multiplier16by16to32_start,_q_multiplier16by16to32_start;
reg  [15:0] _d_doperations2_operand1h,_q_doperations2_operand1h;
reg  [15:0] _d_doperations2_operand1l,_q_doperations2_operand1l;
reg  [15:0] _d_doperations2_operand2h,_q_doperations2_operand2h;
reg  [15:0] _d_doperations2_operand2l,_q_doperations2_operand2l;
reg  [15:0] _d_doperations1_operand1h,_q_doperations1_operand1h;
reg  [15:0] _d_doperations1_operand1l,_q_doperations1_operand1l;
reg  [1:0] _d_index,_q_index;
reg  _p1hz_run;
reg  _timer1hz_run;
reg  _sleepTimer_run;
reg  _timer1khz_run;
reg  _rng_run;
reg  _usend_run;
reg  _background_generator_run;
reg  _tile_map_run;
reg  _bitmap_window_run;
reg  _pixel_writer_run;
reg  _lower_sprites_run;
reg  _upper_sprites_run;
reg  _character_map_window_run;
reg  _terminal_window_run;
reg  _display_run;
reg  _apu_processor_L_run;
reg  _apu_processor_R_run;
reg  _gpu_processor_run;
reg  _divmod32by16to16qr_run;
reg  _divmod16by16to16qr_run;
reg  _multiplier16by16to32_run;
reg  _doperations2_run;
reg  _doperations1_run;
assign out_leds = _q_leds;
assign out_uart_tx = _w_usend_uart_tx;
assign out_audio_l = _w_apu_processor_L_audio_output;
assign out_audio_r = _w_apu_processor_R_audio_output;
assign out_video_r = _w_display_pix_red;
assign out_video_g = _w_display_pix_green;
assign out_video_b = _w_display_pix_blue;
assign out_readData = _d_readData;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_uo_data_in <= 0;
_q_uo_data_in_ready <= 0;
_q_uartInBuffer_addr0 <= 0;
_q_uartInBuffer_wenable1 <= 0;
_q_uartInBuffer_wdata1 <= 0;
_q_uartInBuffer_addr1 <= 0;
_q_uartInBufferNext <= 0;
_q_uartInBufferTop <= 0;
_q_uartOutBuffer_addr0 <= 0;
_q_uartOutBuffer_wenable1 <= 0;
_q_uartOutBuffer_wdata1 <= 0;
_q_uartOutBuffer_addr1 <= 0;
_q_uartOutBufferNext <= 0;
_q_uartOutBufferTop <= 0;
_q_newuartOutBufferTop <= 0;
_q_coProReset <= 0;
_q_delayed_4582_4 <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_uo_data_in <= _d_uo_data_in;
_q_uo_data_in_ready <= _d_uo_data_in_ready;
_q_uartInBuffer_addr0 <= _d_uartInBuffer_addr0;
_q_uartInBuffer_wenable1 <= _d_uartInBuffer_wenable1;
_q_uartInBuffer_wdata1 <= _d_uartInBuffer_wdata1;
_q_uartInBuffer_addr1 <= _d_uartInBuffer_addr1;
_q_uartInBufferNext <= _d_uartInBufferNext;
_q_uartInBufferTop <= _d_uartInBufferTop;
_q_uartOutBuffer_addr0 <= _d_uartOutBuffer_addr0;
_q_uartOutBuffer_wenable1 <= _d_uartOutBuffer_wenable1;
_q_uartOutBuffer_wdata1 <= _d_uartOutBuffer_wdata1;
_q_uartOutBuffer_addr1 <= _d_uartOutBuffer_addr1;
_q_uartOutBufferNext <= _d_uartOutBufferNext;
_q_uartOutBufferTop <= _d_uartOutBufferTop;
_q_newuartOutBufferTop <= _d_newuartOutBufferTop;
_q_coProReset <= _d_coProReset;
_q_delayed_4582_4 <= _d_delayed_4582_4;
_q_leds <= _d_leds;
_q_readData <= _d_readData;
_q_index <= _d_index;
  end
_q_p1hz_resetCounter <= _d_p1hz_resetCounter;
_q_timer1hz_resetCounter <= _d_timer1hz_resetCounter;
_q_sleepTimer_resetCount <= _d_sleepTimer_resetCount;
_q_sleepTimer_resetCounter <= _d_sleepTimer_resetCounter;
_q_timer1khz_resetCount <= _d_timer1khz_resetCount;
_q_timer1khz_resetCounter <= _d_timer1khz_resetCounter;
_q_rng_resetRandom <= _d_rng_resetRandom;
_q_background_generator_backgroundcolour <= _d_background_generator_backgroundcolour;
_q_background_generator_backgroundcolour_alt <= _d_background_generator_backgroundcolour_alt;
_q_background_generator_backgroundcolour_mode <= _d_background_generator_backgroundcolour_mode;
_q_background_generator_background_write <= _d_background_generator_background_write;
_q_tile_map_tm_x <= _d_tile_map_tm_x;
_q_tile_map_tm_y <= _d_tile_map_tm_y;
_q_tile_map_tm_character <= _d_tile_map_tm_character;
_q_tile_map_tm_foreground <= _d_tile_map_tm_foreground;
_q_tile_map_tm_background <= _d_tile_map_tm_background;
_q_tile_map_tm_write <= _d_tile_map_tm_write;
_q_tile_map_tile_writer_tile <= _d_tile_map_tile_writer_tile;
_q_tile_map_tile_writer_line <= _d_tile_map_tile_writer_line;
_q_tile_map_tile_writer_bitmap <= _d_tile_map_tile_writer_bitmap;
_q_tile_map_tm_scrollwrap <= _d_tile_map_tm_scrollwrap;
_q_bitmap_window_bitmap_write_offset <= _d_bitmap_window_bitmap_write_offset;
_q_bitmap_window_bitmap_x_read <= _d_bitmap_window_bitmap_x_read;
_q_bitmap_window_bitmap_y_read <= _d_bitmap_window_bitmap_y_read;
_q_lower_sprites_sprite_set_number <= _d_lower_sprites_sprite_set_number;
_q_lower_sprites_sprite_set_active <= _d_lower_sprites_sprite_set_active;
_q_lower_sprites_sprite_set_double <= _d_lower_sprites_sprite_set_double;
_q_lower_sprites_sprite_set_colour <= _d_lower_sprites_sprite_set_colour;
_q_lower_sprites_sprite_set_x <= _d_lower_sprites_sprite_set_x;
_q_lower_sprites_sprite_set_y <= _d_lower_sprites_sprite_set_y;
_q_lower_sprites_sprite_set_tile <= _d_lower_sprites_sprite_set_tile;
_q_lower_sprites_sprite_layer_write <= _d_lower_sprites_sprite_layer_write;
_q_lower_sprites_sprite_update <= _d_lower_sprites_sprite_update;
_q_lower_sprites_sprite_writer_sprite <= _d_lower_sprites_sprite_writer_sprite;
_q_lower_sprites_sprite_writer_line <= _d_lower_sprites_sprite_writer_line;
_q_lower_sprites_sprite_writer_bitmap <= _d_lower_sprites_sprite_writer_bitmap;
_q_lower_sprites_sprite_writer_active <= _d_lower_sprites_sprite_writer_active;
_q_upper_sprites_sprite_set_number <= _d_upper_sprites_sprite_set_number;
_q_upper_sprites_sprite_set_active <= _d_upper_sprites_sprite_set_active;
_q_upper_sprites_sprite_set_double <= _d_upper_sprites_sprite_set_double;
_q_upper_sprites_sprite_set_colour <= _d_upper_sprites_sprite_set_colour;
_q_upper_sprites_sprite_set_x <= _d_upper_sprites_sprite_set_x;
_q_upper_sprites_sprite_set_y <= _d_upper_sprites_sprite_set_y;
_q_upper_sprites_sprite_set_tile <= _d_upper_sprites_sprite_set_tile;
_q_upper_sprites_sprite_layer_write <= _d_upper_sprites_sprite_layer_write;
_q_upper_sprites_sprite_update <= _d_upper_sprites_sprite_update;
_q_upper_sprites_sprite_writer_sprite <= _d_upper_sprites_sprite_writer_sprite;
_q_upper_sprites_sprite_writer_line <= _d_upper_sprites_sprite_writer_line;
_q_upper_sprites_sprite_writer_bitmap <= _d_upper_sprites_sprite_writer_bitmap;
_q_upper_sprites_sprite_writer_active <= _d_upper_sprites_sprite_writer_active;
_q_character_map_window_tpu_x <= _d_character_map_window_tpu_x;
_q_character_map_window_tpu_y <= _d_character_map_window_tpu_y;
_q_character_map_window_tpu_character <= _d_character_map_window_tpu_character;
_q_character_map_window_tpu_foreground <= _d_character_map_window_tpu_foreground;
_q_character_map_window_tpu_background <= _d_character_map_window_tpu_background;
_q_character_map_window_tpu_write <= _d_character_map_window_tpu_write;
_q_terminal_window_terminal_character <= _d_terminal_window_terminal_character;
_q_terminal_window_terminal_write <= _d_terminal_window_terminal_write;
_q_terminal_window_showterminal <= _d_terminal_window_showterminal;
_q_apu_processor_L_waveform <= _d_apu_processor_L_waveform;
_q_apu_processor_L_note <= _d_apu_processor_L_note;
_q_apu_processor_L_duration <= _d_apu_processor_L_duration;
_q_apu_processor_L_apu_write <= _d_apu_processor_L_apu_write;
_q_apu_processor_R_waveform <= _d_apu_processor_R_waveform;
_q_apu_processor_R_note <= _d_apu_processor_R_note;
_q_apu_processor_R_duration <= _d_apu_processor_R_duration;
_q_apu_processor_R_apu_write <= _d_apu_processor_R_apu_write;
_q_gpu_processor_gpu_x <= _d_gpu_processor_gpu_x;
_q_gpu_processor_gpu_y <= _d_gpu_processor_gpu_y;
_q_gpu_processor_gpu_colour <= _d_gpu_processor_gpu_colour;
_q_gpu_processor_gpu_param0 <= _d_gpu_processor_gpu_param0;
_q_gpu_processor_gpu_param1 <= _d_gpu_processor_gpu_param1;
_q_gpu_processor_gpu_param2 <= _d_gpu_processor_gpu_param2;
_q_gpu_processor_gpu_param3 <= _d_gpu_processor_gpu_param3;
_q_gpu_processor_gpu_write <= _d_gpu_processor_gpu_write;
_q_gpu_processor_blit1_writer_tile <= _d_gpu_processor_blit1_writer_tile;
_q_gpu_processor_blit1_writer_line <= _d_gpu_processor_blit1_writer_line;
_q_gpu_processor_blit1_writer_bitmap <= _d_gpu_processor_blit1_writer_bitmap;
_q_gpu_processor_vector_block_number <= _d_gpu_processor_vector_block_number;
_q_gpu_processor_vector_block_colour <= _d_gpu_processor_vector_block_colour;
_q_gpu_processor_vector_block_xc <= _d_gpu_processor_vector_block_xc;
_q_gpu_processor_vector_block_yc <= _d_gpu_processor_vector_block_yc;
_q_gpu_processor_draw_vector <= _d_gpu_processor_draw_vector;
_q_gpu_processor_vertices_writer_block <= _d_gpu_processor_vertices_writer_block;
_q_gpu_processor_vertices_writer_vertex <= _d_gpu_processor_vertices_writer_vertex;
_q_gpu_processor_vertices_writer_xdelta <= _d_gpu_processor_vertices_writer_xdelta;
_q_gpu_processor_vertices_writer_ydelta <= _d_gpu_processor_vertices_writer_ydelta;
_q_gpu_processor_vertices_writer_active <= _d_gpu_processor_vertices_writer_active;
_q_divmod32by16to16qr_dividendh <= _d_divmod32by16to16qr_dividendh;
_q_divmod32by16to16qr_dividendl <= _d_divmod32by16to16qr_dividendl;
_q_divmod32by16to16qr_divisor <= _d_divmod32by16to16qr_divisor;
_q_divmod32by16to16qr_start <= _d_divmod32by16to16qr_start;
_q_divmod16by16to16qr_dividend <= _d_divmod16by16to16qr_dividend;
_q_divmod16by16to16qr_divisor <= _d_divmod16by16to16qr_divisor;
_q_divmod16by16to16qr_start <= _d_divmod16by16to16qr_start;
_q_multiplier16by16to32_factor1 <= _d_multiplier16by16to32_factor1;
_q_multiplier16by16to32_factor2 <= _d_multiplier16by16to32_factor2;
_q_multiplier16by16to32_start <= _d_multiplier16by16to32_start;
_q_doperations2_operand1h <= _d_doperations2_operand1h;
_q_doperations2_operand1l <= _d_doperations2_operand1l;
_q_doperations2_operand2h <= _d_doperations2_operand2h;
_q_doperations2_operand2l <= _d_doperations2_operand2l;
_q_doperations1_operand1h <= _d_doperations1_operand1h;
_q_doperations1_operand1l <= _d_doperations1_operand1l;
end

M_pulse1hz p1hz (
.in_resetCounter(_d_p1hz_resetCounter),
.out_counter1hz(_w_p1hz_counter1hz),
.out_done(_w_p1hz_done),
.in_run(_p1hz_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_pulse1hz timer1hz (
.in_resetCounter(_d_timer1hz_resetCounter),
.out_counter1hz(_w_timer1hz_counter1hz),
.out_done(_w_timer1hz_done),
.in_run(_timer1hz_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_pulse1khz sleepTimer (
.in_resetCount(_d_sleepTimer_resetCount),
.in_resetCounter(_d_sleepTimer_resetCounter),
.out_counter1khz(_w_sleepTimer_counter1khz),
.out_done(_w_sleepTimer_done),
.in_run(_sleepTimer_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_pulse1khz timer1khz (
.in_resetCount(_d_timer1khz_resetCount),
.in_resetCounter(_d_timer1khz_resetCounter),
.out_counter1khz(_w_timer1khz_counter1khz),
.out_done(_w_timer1khz_done),
.in_run(_timer1khz_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_random rng (
.in_resetRandom(_d_rng_resetRandom),
.out_g_noise_out(_w_rng_g_noise_out),
.out_u_noise_out(_w_rng_u_noise_out),
.out_done(_w_rng_done),
.in_run(_rng_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_uart_sender #(
.IO_DATA_IN_WIDTH(8),
.IO_DATA_IN_INIT(0),
.IO_DATA_IN_SIGNED(0),
.IO_DATA_IN_READY_WIDTH(1),
.IO_DATA_IN_READY_INIT(0),
.IO_DATA_IN_READY_SIGNED(0),
.IO_BUSY_WIDTH(1),
.IO_BUSY_INIT(0),
.IO_BUSY_SIGNED(0)
) usend (
.in_io_data_in(_d_uo_data_in),
.in_io_data_in_ready(_d_uo_data_in_ready),
.out_io_busy(_w_usend_io_busy),
.out_uart_tx(_w_usend_uart_tx),
.out_done(_w_usend_done),
.in_run(_usend_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_uart_receiver #(
.IO_DATA_OUT_WIDTH(8),
.IO_DATA_OUT_INIT(0),
.IO_DATA_OUT_SIGNED(0),
.IO_DATA_OUT_READY_WIDTH(1),
.IO_DATA_OUT_READY_INIT(0),
.IO_DATA_OUT_READY_SIGNED(0)
) urecv (
.in_uart_rx(in_uart_rx),
.out_io_data_out(_w_urecv_io_data_out),
.out_io_data_out_ready(_w_urecv_io_data_out_ready),
.reset(reset),
.clock(in_clock_50mhz)
);
M_background background_generator (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_staticGenerator(_w_rng_g_noise_out),
.in_backgroundcolour(_d_background_generator_backgroundcolour),
.in_backgroundcolour_alt(_d_background_generator_backgroundcolour_alt),
.in_backgroundcolour_mode(_d_background_generator_backgroundcolour_mode),
.in_background_write(_d_background_generator_background_write),
.out_pix_red(_w_background_generator_pix_red),
.out_pix_green(_w_background_generator_pix_green),
.out_pix_blue(_w_background_generator_pix_blue),
.out_done(_w_background_generator_done),
.in_run(_background_generator_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_tilemap tile_map (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_tm_x(_d_tile_map_tm_x),
.in_tm_y(_d_tile_map_tm_y),
.in_tm_character(_d_tile_map_tm_character),
.in_tm_foreground(_d_tile_map_tm_foreground),
.in_tm_background(_d_tile_map_tm_background),
.in_tm_write(_d_tile_map_tm_write),
.in_tile_writer_tile(_d_tile_map_tile_writer_tile),
.in_tile_writer_line(_d_tile_map_tile_writer_line),
.in_tile_writer_bitmap(_d_tile_map_tile_writer_bitmap),
.in_tm_scrollwrap(_d_tile_map_tm_scrollwrap),
.out_pix_red(_w_tile_map_pix_red),
.out_pix_green(_w_tile_map_pix_green),
.out_pix_blue(_w_tile_map_pix_blue),
.out_tilemap_display(_w_tile_map_tilemap_display),
.out_tm_lastaction(_w_tile_map_tm_lastaction),
.out_tm_active(_w_tile_map_tm_active),
.out_done(_w_tile_map_done),
.in_run(_tile_map_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_bitmap #(
.BITMAP_ADDR0_WIDTH(19),
.BITMAP_ADDR0_INIT(0),
.BITMAP_ADDR0_SIGNED(0),
.BITMAP_RDATA0_WIDTH(7),
.BITMAP_RDATA0_INIT(0),
.BITMAP_RDATA0_SIGNED(0)
) bitmap_window (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_bitmap_write_offset(_d_bitmap_window_bitmap_write_offset),
.in_bitmap_x_read(_d_bitmap_window_bitmap_x_read),
.in_bitmap_y_read(_d_bitmap_window_bitmap_y_read),
.in_bitmap_rdata0(_w_mem_bitmap_rdata0),
.out_pix_red(_w_bitmap_window_pix_red),
.out_pix_green(_w_bitmap_window_pix_green),
.out_pix_blue(_w_bitmap_window_pix_blue),
.out_bitmap_display(_w_bitmap_window_bitmap_display),
.out_x_offset(_w_bitmap_window_x_offset),
.out_y_offset(_w_bitmap_window_y_offset),
.out_bitmap_colour_read(_w_bitmap_window_bitmap_colour_read),
.out_bitmap_addr0(_w_bitmap_window_bitmap_addr0),
.out_done(_w_bitmap_window_done),
.in_run(_bitmap_window_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_bitmapwriter #(
.BITMAP_ADDR1_WIDTH(19),
.BITMAP_ADDR1_INIT(0),
.BITMAP_ADDR1_SIGNED(0),
.BITMAP_WENABLE1_WIDTH(1),
.BITMAP_WENABLE1_INIT(0),
.BITMAP_WENABLE1_SIGNED(0),
.BITMAP_WDATA1_WIDTH(7),
.BITMAP_WDATA1_INIT(0),
.BITMAP_WDATA1_SIGNED(0)
) pixel_writer (
.in_bitmap_x_write(_w_gpu_processor_bitmap_x_write),
.in_bitmap_y_write(_w_gpu_processor_bitmap_y_write),
.in_bitmap_colour_write(_w_gpu_processor_bitmap_colour_write),
.in_bitmap_write(_w_gpu_processor_bitmap_write),
.in_x_offset(_w_bitmap_window_x_offset),
.in_y_offset(_w_bitmap_window_y_offset),
.out_bitmap_addr1(_w_pixel_writer_bitmap_addr1),
.out_bitmap_wenable1(_w_pixel_writer_bitmap_wenable1),
.out_bitmap_wdata1(_w_pixel_writer_bitmap_wdata1),
.out_done(_w_pixel_writer_done),
.in_run(_pixel_writer_run),
.reset(reset),
.clock(in_video_clock)
);
M_sprite_layer lower_sprites (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_sprite_set_number(_d_lower_sprites_sprite_set_number),
.in_sprite_set_active(_d_lower_sprites_sprite_set_active),
.in_sprite_set_double(_d_lower_sprites_sprite_set_double),
.in_sprite_set_colour(_d_lower_sprites_sprite_set_colour),
.in_sprite_set_x(_d_lower_sprites_sprite_set_x),
.in_sprite_set_y(_d_lower_sprites_sprite_set_y),
.in_sprite_set_tile(_d_lower_sprites_sprite_set_tile),
.in_sprite_layer_write(_d_lower_sprites_sprite_layer_write),
.in_sprite_update(_d_lower_sprites_sprite_update),
.in_collision_layer_1(_w_bitmap_window_bitmap_display),
.in_collision_layer_2(_w_tile_map_tilemap_display),
.in_collision_layer_3(_w_upper_sprites_sprite_layer_display),
.in_sprite_writer_sprite(_d_lower_sprites_sprite_writer_sprite),
.in_sprite_writer_line(_d_lower_sprites_sprite_writer_line),
.in_sprite_writer_bitmap(_d_lower_sprites_sprite_writer_bitmap),
.in_sprite_writer_active(_d_lower_sprites_sprite_writer_active),
.out_pix_red(_w_lower_sprites_pix_red),
.out_pix_green(_w_lower_sprites_pix_green),
.out_pix_blue(_w_lower_sprites_pix_blue),
.out_sprite_layer_display(_w_lower_sprites_sprite_layer_display),
.out_sprite_read_active(_w_lower_sprites_sprite_read_active),
.out_sprite_read_double(_w_lower_sprites_sprite_read_double),
.out_sprite_read_colour(_w_lower_sprites_sprite_read_colour),
.out_sprite_read_x(_w_lower_sprites_sprite_read_x),
.out_sprite_read_y(_w_lower_sprites_sprite_read_y),
.out_sprite_read_tile(_w_lower_sprites_sprite_read_tile),
.out_collision_0(_w_lower_sprites_collision_0),
.out_collision_1(_w_lower_sprites_collision_1),
.out_collision_2(_w_lower_sprites_collision_2),
.out_collision_3(_w_lower_sprites_collision_3),
.out_collision_4(_w_lower_sprites_collision_4),
.out_collision_5(_w_lower_sprites_collision_5),
.out_collision_6(_w_lower_sprites_collision_6),
.out_collision_7(_w_lower_sprites_collision_7),
.out_collision_8(_w_lower_sprites_collision_8),
.out_collision_9(_w_lower_sprites_collision_9),
.out_collision_10(_w_lower_sprites_collision_10),
.out_collision_11(_w_lower_sprites_collision_11),
.out_collision_12(_w_lower_sprites_collision_12),
.out_done(_w_lower_sprites_done),
.in_run(_lower_sprites_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_sprite_layer upper_sprites (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_sprite_set_number(_d_upper_sprites_sprite_set_number),
.in_sprite_set_active(_d_upper_sprites_sprite_set_active),
.in_sprite_set_double(_d_upper_sprites_sprite_set_double),
.in_sprite_set_colour(_d_upper_sprites_sprite_set_colour),
.in_sprite_set_x(_d_upper_sprites_sprite_set_x),
.in_sprite_set_y(_d_upper_sprites_sprite_set_y),
.in_sprite_set_tile(_d_upper_sprites_sprite_set_tile),
.in_sprite_layer_write(_d_upper_sprites_sprite_layer_write),
.in_sprite_update(_d_upper_sprites_sprite_update),
.in_collision_layer_1(_w_bitmap_window_bitmap_display),
.in_collision_layer_2(_w_tile_map_tilemap_display),
.in_collision_layer_3(_w_lower_sprites_sprite_layer_display),
.in_sprite_writer_sprite(_d_upper_sprites_sprite_writer_sprite),
.in_sprite_writer_line(_d_upper_sprites_sprite_writer_line),
.in_sprite_writer_bitmap(_d_upper_sprites_sprite_writer_bitmap),
.in_sprite_writer_active(_d_upper_sprites_sprite_writer_active),
.out_pix_red(_w_upper_sprites_pix_red),
.out_pix_green(_w_upper_sprites_pix_green),
.out_pix_blue(_w_upper_sprites_pix_blue),
.out_sprite_layer_display(_w_upper_sprites_sprite_layer_display),
.out_sprite_read_active(_w_upper_sprites_sprite_read_active),
.out_sprite_read_double(_w_upper_sprites_sprite_read_double),
.out_sprite_read_colour(_w_upper_sprites_sprite_read_colour),
.out_sprite_read_x(_w_upper_sprites_sprite_read_x),
.out_sprite_read_y(_w_upper_sprites_sprite_read_y),
.out_sprite_read_tile(_w_upper_sprites_sprite_read_tile),
.out_collision_0(_w_upper_sprites_collision_0),
.out_collision_1(_w_upper_sprites_collision_1),
.out_collision_2(_w_upper_sprites_collision_2),
.out_collision_3(_w_upper_sprites_collision_3),
.out_collision_4(_w_upper_sprites_collision_4),
.out_collision_5(_w_upper_sprites_collision_5),
.out_collision_6(_w_upper_sprites_collision_6),
.out_collision_7(_w_upper_sprites_collision_7),
.out_collision_8(_w_upper_sprites_collision_8),
.out_collision_9(_w_upper_sprites_collision_9),
.out_collision_10(_w_upper_sprites_collision_10),
.out_collision_11(_w_upper_sprites_collision_11),
.out_collision_12(_w_upper_sprites_collision_12),
.out_done(_w_upper_sprites_done),
.in_run(_upper_sprites_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_character_map character_map_window (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_tpu_x(_d_character_map_window_tpu_x),
.in_tpu_y(_d_character_map_window_tpu_y),
.in_tpu_character(_d_character_map_window_tpu_character),
.in_tpu_foreground(_d_character_map_window_tpu_foreground),
.in_tpu_background(_d_character_map_window_tpu_background),
.in_tpu_write(_d_character_map_window_tpu_write),
.out_pix_red(_w_character_map_window_pix_red),
.out_pix_green(_w_character_map_window_pix_green),
.out_pix_blue(_w_character_map_window_pix_blue),
.out_character_map_display(_w_character_map_window_character_map_display),
.out_tpu_active(_w_character_map_window_tpu_active),
.out_done(_w_character_map_window_done),
.in_run(_character_map_window_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_terminal terminal_window (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_terminal_character(_d_terminal_window_terminal_character),
.in_terminal_write(_d_terminal_window_terminal_write),
.in_showterminal(_d_terminal_window_showterminal),
.in_timer1hz(_w_p1hz_counter1hz),
.out_pix_red(_w_terminal_window_pix_red),
.out_pix_green(_w_terminal_window_pix_green),
.out_pix_blue(_w_terminal_window_pix_blue),
.out_terminal_display(_w_terminal_window_terminal_display),
.out_terminal_active(_w_terminal_window_terminal_active),
.out_done(_w_terminal_window_done),
.in_run(_terminal_window_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_multiplex_display display (
.in_pix_x(in_pix_x),
.in_pix_y(in_pix_y),
.in_pix_active(in_pix_active),
.in_pix_vblank(in_vblank),
.in_background_r(_w_background_generator_pix_red),
.in_background_g(_w_background_generator_pix_green),
.in_background_b(_w_background_generator_pix_blue),
.in_tilemap_r(_w_tile_map_pix_red),
.in_tilemap_g(_w_tile_map_pix_green),
.in_tilemap_b(_w_tile_map_pix_blue),
.in_tilemap_display(_w_tile_map_tilemap_display),
.in_lower_sprites_r(_w_lower_sprites_pix_red),
.in_lower_sprites_g(_w_lower_sprites_pix_green),
.in_lower_sprites_b(_w_lower_sprites_pix_blue),
.in_lower_sprites_display(_w_lower_sprites_sprite_layer_display),
.in_bitmap_r(_w_bitmap_window_pix_red),
.in_bitmap_g(_w_bitmap_window_pix_green),
.in_bitmap_b(_w_bitmap_window_pix_blue),
.in_bitmap_display(_w_bitmap_window_bitmap_display),
.in_upper_sprites_r(_w_upper_sprites_pix_red),
.in_upper_sprites_g(_w_upper_sprites_pix_green),
.in_upper_sprites_b(_w_upper_sprites_pix_blue),
.in_upper_sprites_display(_w_upper_sprites_sprite_layer_display),
.in_character_map_r(_w_character_map_window_pix_red),
.in_character_map_g(_w_character_map_window_pix_green),
.in_character_map_b(_w_character_map_window_pix_blue),
.in_character_map_display(_w_character_map_window_character_map_display),
.in_terminal_r(_w_terminal_window_pix_red),
.in_terminal_g(_w_terminal_window_pix_green),
.in_terminal_b(_w_terminal_window_pix_blue),
.in_terminal_display(_w_terminal_window_terminal_display),
.out_pix_red(_w_display_pix_red),
.out_pix_green(_w_display_pix_green),
.out_pix_blue(_w_display_pix_blue),
.out_done(_w_display_done),
.in_run(_display_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_apu apu_processor_L (
.in_waveform(_d_apu_processor_L_waveform),
.in_note(_d_apu_processor_L_note),
.in_duration(_d_apu_processor_L_duration),
.in_apu_write(_d_apu_processor_L_apu_write),
.in_staticGenerator(_w_rng_g_noise_out),
.out_audio_active(_w_apu_processor_L_audio_active),
.out_audio_output(_w_apu_processor_L_audio_output),
.out_done(_w_apu_processor_L_done),
.in_run(_apu_processor_L_run),
.reset(reset),
.clock(in_clock_25mhz)
);
M_apu apu_processor_R (
.in_waveform(_d_apu_processor_R_waveform),
.in_note(_d_apu_processor_R_note),
.in_duration(_d_apu_processor_R_duration),
.in_apu_write(_d_apu_processor_R_apu_write),
.in_staticGenerator(_w_rng_g_noise_out),
.out_audio_active(_w_apu_processor_R_audio_active),
.out_audio_output(_w_apu_processor_R_audio_output),
.out_done(_w_apu_processor_R_done),
.in_run(_apu_processor_R_run),
.reset(reset),
.clock(in_clock_25mhz)
);
M_gpu gpu_processor (
.in_gpu_x(_d_gpu_processor_gpu_x),
.in_gpu_y(_d_gpu_processor_gpu_y),
.in_gpu_colour(_d_gpu_processor_gpu_colour),
.in_gpu_param0(_d_gpu_processor_gpu_param0),
.in_gpu_param1(_d_gpu_processor_gpu_param1),
.in_gpu_param2(_d_gpu_processor_gpu_param2),
.in_gpu_param3(_d_gpu_processor_gpu_param3),
.in_gpu_write(_d_gpu_processor_gpu_write),
.in_blit1_writer_tile(_d_gpu_processor_blit1_writer_tile),
.in_blit1_writer_line(_d_gpu_processor_blit1_writer_line),
.in_blit1_writer_bitmap(_d_gpu_processor_blit1_writer_bitmap),
.in_vector_block_number(_d_gpu_processor_vector_block_number),
.in_vector_block_colour(_d_gpu_processor_vector_block_colour),
.in_vector_block_xc(_d_gpu_processor_vector_block_xc),
.in_vector_block_yc(_d_gpu_processor_vector_block_yc),
.in_draw_vector(_d_gpu_processor_draw_vector),
.in_vertices_writer_block(_d_gpu_processor_vertices_writer_block),
.in_vertices_writer_vertex(_d_gpu_processor_vertices_writer_vertex),
.in_vertices_writer_xdelta(_d_gpu_processor_vertices_writer_xdelta),
.in_vertices_writer_ydelta(_d_gpu_processor_vertices_writer_ydelta),
.in_vertices_writer_active(_d_gpu_processor_vertices_writer_active),
.out_bitmap_x_write(_w_gpu_processor_bitmap_x_write),
.out_bitmap_y_write(_w_gpu_processor_bitmap_y_write),
.out_bitmap_colour_write(_w_gpu_processor_bitmap_colour_write),
.out_bitmap_write(_w_gpu_processor_bitmap_write),
.out_gpu_active(_w_gpu_processor_gpu_active),
.out_vector_block_active(_w_gpu_processor_vector_block_active),
.out_done(_w_gpu_processor_done),
.in_run(_gpu_processor_run),
.reset(in_video_reset),
.clock(in_video_clock)
);
M_divmod32by16 divmod32by16to16qr (
.in_dividendh(_d_divmod32by16to16qr_dividendh),
.in_dividendl(_d_divmod32by16to16qr_dividendl),
.in_divisor(_d_divmod32by16to16qr_divisor),
.in_start(_d_divmod32by16to16qr_start),
.out_quotient(_w_divmod32by16to16qr_quotient),
.out_remainder(_w_divmod32by16to16qr_remainder),
.out_active(_w_divmod32by16to16qr_active),
.out_done(_w_divmod32by16to16qr_done),
.in_run(_divmod32by16to16qr_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_divmod16by16 divmod16by16to16qr (
.in_dividend(_d_divmod16by16to16qr_dividend),
.in_divisor(_d_divmod16by16to16qr_divisor),
.in_start(_d_divmod16by16to16qr_start),
.out_quotient(_w_divmod16by16to16qr_quotient),
.out_remainder(_w_divmod16by16to16qr_remainder),
.out_active(_w_divmod16by16to16qr_active),
.out_done(_w_divmod16by16to16qr_done),
.in_run(_divmod16by16to16qr_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_multi16by16to32DSP multiplier16by16to32 (
.in_factor1(_d_multiplier16by16to32_factor1),
.in_factor2(_d_multiplier16by16to32_factor2),
.in_start(_d_multiplier16by16to32_start),
.out_product(_w_multiplier16by16to32_product),
.out_active(_w_multiplier16by16to32_active),
.out_done(_w_multiplier16by16to32_done),
.in_run(_multiplier16by16to32_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_doubleaddsub2input doperations2 (
.in_operand1h(_d_doperations2_operand1h),
.in_operand1l(_d_doperations2_operand1l),
.in_operand2h(_d_doperations2_operand2h),
.in_operand2l(_d_doperations2_operand2l),
.out_total(_w_doperations2_total),
.out_difference(_w_doperations2_difference),
.out_binaryxor(_w_doperations2_binaryxor),
.out_binaryor(_w_doperations2_binaryor),
.out_binaryand(_w_doperations2_binaryand),
.out_maximum(_w_doperations2_maximum),
.out_minimum(_w_doperations2_minimum),
.out_equal(_w_doperations2_equal),
.out_lessthan(_w_doperations2_lessthan),
.out_done(_w_doperations2_done),
.in_run(_doperations2_run),
.reset(reset),
.clock(in_clock_50mhz)
);
M_doubleaddsub1input doperations1 (
.in_operand1h(_d_doperations1_operand1h),
.in_operand1l(_d_doperations1_operand1l),
.out_increment(_w_doperations1_increment),
.out_decrement(_w_doperations1_decrement),
.out_times2(_w_doperations1_times2),
.out_divide2(_w_doperations1_divide2),
.out_negation(_w_doperations1_negation),
.out_binaryinvert(_w_doperations1_binaryinvert),
.out_absolute(_w_doperations1_absolute),
.out_zeroequal(_w_doperations1_zeroequal),
.out_zeroless(_w_doperations1_zeroless),
.out_done(_w_doperations1_done),
.in_run(_doperations1_run),
.reset(reset),
.clock(in_clock_50mhz)
);

M_memmap_io_mem_bitmap __mem__bitmap(
.clock0(in_video_clock),
.clock1(in_video_clock),
.in_bitmap_addr0(_w_bitmap_window_bitmap_addr0),
.in_bitmap_wenable1(_w_pixel_writer_bitmap_wenable1),
.in_bitmap_wdata1(_w_pixel_writer_bitmap_wdata1),
.in_bitmap_addr1(_w_pixel_writer_bitmap_addr1),
.out_bitmap_rdata0(_w_mem_bitmap_rdata0)
);
M_memmap_io_mem_uartInBuffer __mem__uartInBuffer(
.clock0(clock),
.clock1(clock),
.in_uartInBuffer_addr0(_d_uartInBuffer_addr0),
.in_uartInBuffer_wenable1(_d_uartInBuffer_wenable1),
.in_uartInBuffer_wdata1(_d_uartInBuffer_wdata1),
.in_uartInBuffer_addr1(_d_uartInBuffer_addr1),
.out_uartInBuffer_rdata0(_w_mem_uartInBuffer_rdata0)
);
M_memmap_io_mem_uartOutBuffer __mem__uartOutBuffer(
.clock0(clock),
.clock1(clock),
.in_uartOutBuffer_addr0(_d_uartOutBuffer_addr0),
.in_uartOutBuffer_wenable1(_d_uartOutBuffer_wenable1),
.in_uartOutBuffer_wdata1(_d_uartOutBuffer_wdata1),
.in_uartOutBuffer_addr1(_d_uartOutBuffer_addr1),
.out_uartOutBuffer_rdata0(_w_mem_uartOutBuffer_rdata0)
);


always @* begin
_d_uo_data_in = _q_uo_data_in;
_d_uo_data_in_ready = _q_uo_data_in_ready;
_d_uartInBuffer_addr0 = _q_uartInBuffer_addr0;
_d_uartInBuffer_wenable1 = _q_uartInBuffer_wenable1;
_d_uartInBuffer_wdata1 = _q_uartInBuffer_wdata1;
_d_uartInBuffer_addr1 = _q_uartInBuffer_addr1;
_d_uartInBufferNext = _q_uartInBufferNext;
_d_uartInBufferTop = _q_uartInBufferTop;
_d_uartOutBuffer_addr0 = _q_uartOutBuffer_addr0;
_d_uartOutBuffer_wenable1 = _q_uartOutBuffer_wenable1;
_d_uartOutBuffer_wdata1 = _q_uartOutBuffer_wdata1;
_d_uartOutBuffer_addr1 = _q_uartOutBuffer_addr1;
_d_uartOutBufferNext = _q_uartOutBufferNext;
_d_uartOutBufferTop = _q_uartOutBufferTop;
_d_newuartOutBufferTop = _q_newuartOutBufferTop;
_d_coProReset = _q_coProReset;
_d_delayed_4582_4 = _q_delayed_4582_4;
_d_leds = _q_leds;
_d_readData = _q_readData;
_d_p1hz_resetCounter = _q_p1hz_resetCounter;
_d_timer1hz_resetCounter = _q_timer1hz_resetCounter;
_d_sleepTimer_resetCount = _q_sleepTimer_resetCount;
_d_sleepTimer_resetCounter = _q_sleepTimer_resetCounter;
_d_timer1khz_resetCount = _q_timer1khz_resetCount;
_d_timer1khz_resetCounter = _q_timer1khz_resetCounter;
_d_rng_resetRandom = _q_rng_resetRandom;
_d_background_generator_backgroundcolour = _q_background_generator_backgroundcolour;
_d_background_generator_backgroundcolour_alt = _q_background_generator_backgroundcolour_alt;
_d_background_generator_backgroundcolour_mode = _q_background_generator_backgroundcolour_mode;
_d_background_generator_background_write = _q_background_generator_background_write;
_d_tile_map_tm_x = _q_tile_map_tm_x;
_d_tile_map_tm_y = _q_tile_map_tm_y;
_d_tile_map_tm_character = _q_tile_map_tm_character;
_d_tile_map_tm_foreground = _q_tile_map_tm_foreground;
_d_tile_map_tm_background = _q_tile_map_tm_background;
_d_tile_map_tm_write = _q_tile_map_tm_write;
_d_tile_map_tile_writer_tile = _q_tile_map_tile_writer_tile;
_d_tile_map_tile_writer_line = _q_tile_map_tile_writer_line;
_d_tile_map_tile_writer_bitmap = _q_tile_map_tile_writer_bitmap;
_d_tile_map_tm_scrollwrap = _q_tile_map_tm_scrollwrap;
_d_bitmap_window_bitmap_write_offset = _q_bitmap_window_bitmap_write_offset;
_d_bitmap_window_bitmap_x_read = _q_bitmap_window_bitmap_x_read;
_d_bitmap_window_bitmap_y_read = _q_bitmap_window_bitmap_y_read;
_d_lower_sprites_sprite_set_number = _q_lower_sprites_sprite_set_number;
_d_lower_sprites_sprite_set_active = _q_lower_sprites_sprite_set_active;
_d_lower_sprites_sprite_set_double = _q_lower_sprites_sprite_set_double;
_d_lower_sprites_sprite_set_colour = _q_lower_sprites_sprite_set_colour;
_d_lower_sprites_sprite_set_x = _q_lower_sprites_sprite_set_x;
_d_lower_sprites_sprite_set_y = _q_lower_sprites_sprite_set_y;
_d_lower_sprites_sprite_set_tile = _q_lower_sprites_sprite_set_tile;
_d_lower_sprites_sprite_layer_write = _q_lower_sprites_sprite_layer_write;
_d_lower_sprites_sprite_update = _q_lower_sprites_sprite_update;
_d_lower_sprites_sprite_writer_sprite = _q_lower_sprites_sprite_writer_sprite;
_d_lower_sprites_sprite_writer_line = _q_lower_sprites_sprite_writer_line;
_d_lower_sprites_sprite_writer_bitmap = _q_lower_sprites_sprite_writer_bitmap;
_d_lower_sprites_sprite_writer_active = _q_lower_sprites_sprite_writer_active;
_d_upper_sprites_sprite_set_number = _q_upper_sprites_sprite_set_number;
_d_upper_sprites_sprite_set_active = _q_upper_sprites_sprite_set_active;
_d_upper_sprites_sprite_set_double = _q_upper_sprites_sprite_set_double;
_d_upper_sprites_sprite_set_colour = _q_upper_sprites_sprite_set_colour;
_d_upper_sprites_sprite_set_x = _q_upper_sprites_sprite_set_x;
_d_upper_sprites_sprite_set_y = _q_upper_sprites_sprite_set_y;
_d_upper_sprites_sprite_set_tile = _q_upper_sprites_sprite_set_tile;
_d_upper_sprites_sprite_layer_write = _q_upper_sprites_sprite_layer_write;
_d_upper_sprites_sprite_update = _q_upper_sprites_sprite_update;
_d_upper_sprites_sprite_writer_sprite = _q_upper_sprites_sprite_writer_sprite;
_d_upper_sprites_sprite_writer_line = _q_upper_sprites_sprite_writer_line;
_d_upper_sprites_sprite_writer_bitmap = _q_upper_sprites_sprite_writer_bitmap;
_d_upper_sprites_sprite_writer_active = _q_upper_sprites_sprite_writer_active;
_d_character_map_window_tpu_x = _q_character_map_window_tpu_x;
_d_character_map_window_tpu_y = _q_character_map_window_tpu_y;
_d_character_map_window_tpu_character = _q_character_map_window_tpu_character;
_d_character_map_window_tpu_foreground = _q_character_map_window_tpu_foreground;
_d_character_map_window_tpu_background = _q_character_map_window_tpu_background;
_d_character_map_window_tpu_write = _q_character_map_window_tpu_write;
_d_terminal_window_terminal_character = _q_terminal_window_terminal_character;
_d_terminal_window_terminal_write = _q_terminal_window_terminal_write;
_d_terminal_window_showterminal = _q_terminal_window_showterminal;
_d_apu_processor_L_waveform = _q_apu_processor_L_waveform;
_d_apu_processor_L_note = _q_apu_processor_L_note;
_d_apu_processor_L_duration = _q_apu_processor_L_duration;
_d_apu_processor_L_apu_write = _q_apu_processor_L_apu_write;
_d_apu_processor_R_waveform = _q_apu_processor_R_waveform;
_d_apu_processor_R_note = _q_apu_processor_R_note;
_d_apu_processor_R_duration = _q_apu_processor_R_duration;
_d_apu_processor_R_apu_write = _q_apu_processor_R_apu_write;
_d_gpu_processor_gpu_x = _q_gpu_processor_gpu_x;
_d_gpu_processor_gpu_y = _q_gpu_processor_gpu_y;
_d_gpu_processor_gpu_colour = _q_gpu_processor_gpu_colour;
_d_gpu_processor_gpu_param0 = _q_gpu_processor_gpu_param0;
_d_gpu_processor_gpu_param1 = _q_gpu_processor_gpu_param1;
_d_gpu_processor_gpu_param2 = _q_gpu_processor_gpu_param2;
_d_gpu_processor_gpu_param3 = _q_gpu_processor_gpu_param3;
_d_gpu_processor_gpu_write = _q_gpu_processor_gpu_write;
_d_gpu_processor_blit1_writer_tile = _q_gpu_processor_blit1_writer_tile;
_d_gpu_processor_blit1_writer_line = _q_gpu_processor_blit1_writer_line;
_d_gpu_processor_blit1_writer_bitmap = _q_gpu_processor_blit1_writer_bitmap;
_d_gpu_processor_vector_block_number = _q_gpu_processor_vector_block_number;
_d_gpu_processor_vector_block_colour = _q_gpu_processor_vector_block_colour;
_d_gpu_processor_vector_block_xc = _q_gpu_processor_vector_block_xc;
_d_gpu_processor_vector_block_yc = _q_gpu_processor_vector_block_yc;
_d_gpu_processor_draw_vector = _q_gpu_processor_draw_vector;
_d_gpu_processor_vertices_writer_block = _q_gpu_processor_vertices_writer_block;
_d_gpu_processor_vertices_writer_vertex = _q_gpu_processor_vertices_writer_vertex;
_d_gpu_processor_vertices_writer_xdelta = _q_gpu_processor_vertices_writer_xdelta;
_d_gpu_processor_vertices_writer_ydelta = _q_gpu_processor_vertices_writer_ydelta;
_d_gpu_processor_vertices_writer_active = _q_gpu_processor_vertices_writer_active;
_d_divmod32by16to16qr_dividendh = _q_divmod32by16to16qr_dividendh;
_d_divmod32by16to16qr_dividendl = _q_divmod32by16to16qr_dividendl;
_d_divmod32by16to16qr_divisor = _q_divmod32by16to16qr_divisor;
_d_divmod32by16to16qr_start = _q_divmod32by16to16qr_start;
_d_divmod16by16to16qr_dividend = _q_divmod16by16to16qr_dividend;
_d_divmod16by16to16qr_divisor = _q_divmod16by16to16qr_divisor;
_d_divmod16by16to16qr_start = _q_divmod16by16to16qr_start;
_d_multiplier16by16to32_factor1 = _q_multiplier16by16to32_factor1;
_d_multiplier16by16to32_factor2 = _q_multiplier16by16to32_factor2;
_d_multiplier16by16to32_start = _q_multiplier16by16to32_start;
_d_doperations2_operand1h = _q_doperations2_operand1h;
_d_doperations2_operand1l = _q_doperations2_operand1l;
_d_doperations2_operand2h = _q_doperations2_operand2h;
_d_doperations2_operand2l = _q_doperations2_operand2l;
_d_doperations1_operand1h = _q_doperations1_operand1h;
_d_doperations1_operand1l = _q_doperations1_operand1l;
_d_index = _q_index;
_p1hz_run = 1;
_timer1hz_run = 1;
_sleepTimer_run = 1;
_timer1khz_run = 1;
_rng_run = 1;
_usend_run = 1;
_background_generator_run = 1;
_tile_map_run = 1;
_bitmap_window_run = 1;
_pixel_writer_run = 1;
_lower_sprites_run = 1;
_upper_sprites_run = 1;
_character_map_window_run = 1;
_terminal_window_run = 1;
_display_run = 1;
_apu_processor_L_run = 1;
_apu_processor_R_run = 1;
_gpu_processor_run = 1;
_divmod32by16to16qr_run = 1;
_divmod16by16to16qr_run = 1;
_multiplier16by16to32_run = 1;
_doperations2_run = 1;
_doperations1_run = 1;
_t_reg_btns = 0;
// _always_pre
_t_reg_btns = _d_delayed_4582_4;
_d_delayed_4582_4 =  in_btns;
_d_uartInBuffer_wenable1 = 1;
_d_uartInBuffer_addr0 = _q_uartInBufferNext;
_d_uartInBuffer_addr1 = _q_uartInBufferTop;
_d_uartOutBuffer_wenable1 = 1;
_d_uartOutBuffer_addr0 = _q_uartOutBufferNext;
_d_uartOutBuffer_addr1 = _q_uartOutBufferTop;
_d_uo_data_in_ready = 0;
_d_divmod32by16to16qr_start = 0;
_d_divmod16by16to16qr_start = 0;
_d_multiplier16by16to32_start = 0;
_d_p1hz_resetCounter = 0;
_d_sleepTimer_resetCounter = 0;
_d_timer1hz_resetCounter = 0;
_d_timer1khz_resetCounter = 0;
_d_rng_resetRandom = 0;
_d_uartInBuffer_wdata1 = _w_urecv_io_data_out;
_d_uartInBufferTop = (_w_urecv_io_data_out_ready)?_q_uartInBufferTop+1:_q_uartInBufferTop;
_d_uo_data_in = _w_mem_uartOutBuffer_rdata0;
_d_uo_data_in_ready = (_q_uartOutBufferNext!=_q_uartOutBufferTop)&&(!_w_usend_io_busy);
_d_uartOutBufferNext = ((_q_uartOutBufferNext!=_q_uartOutBufferTop)&&(!_w_usend_io_busy))?_q_uartOutBufferNext+1:_q_uartOutBufferNext;
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_uo_data_in = 0;
_d_uo_data_in_ready = 0;
_d_uartInBuffer_addr0 = 0;
_d_uartInBuffer_wenable1 = 0;
_d_uartInBuffer_wdata1 = 0;
_d_uartInBuffer_addr1 = 0;
_d_uartInBufferNext = 0;
_d_uartInBufferTop = 0;
_d_uartOutBuffer_addr0 = 0;
_d_uartOutBuffer_wenable1 = 0;
_d_uartOutBuffer_wdata1 = 0;
_d_uartOutBuffer_addr1 = 0;
_d_uartOutBufferNext = 0;
_d_uartOutBufferTop = 0;
_d_newuartOutBufferTop = 0;
_d_coProReset = 0;
_t_reg_btns = 0;
// --
_d_terminal_window_showterminal = 1;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
_d_uartOutBufferTop = _q_newuartOutBufferTop;
if (in_memoryRead) begin
// __block_5
// __block_7
  case (in_memoryAddress[12+:4])
  4'hf: begin
// __block_9_case
// __block_10
  case (in_memoryAddress[8+:4])
  4'h0: begin
// __block_12_case
// __block_13
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_15_case
// __block_16
_d_readData = {8'b0,_w_mem_uartInBuffer_rdata0};
_d_uartInBufferNext = _q_uartInBufferNext+1;
// __block_17
  end
  4'h1: begin
// __block_18_case
// __block_19
_d_readData = {14'b0,(_d_uartOutBufferTop+1==_d_uartOutBufferNext),(_q_uartInBufferNext!=_d_uartInBufferTop)};
// __block_20
  end
  4'h2: begin
// __block_21_case
// __block_22
_d_readData = _q_leds;
// __block_23
  end
  4'h3: begin
// __block_24_case
// __block_25
_d_readData = {9'b0,_t_reg_btns[0+:7]};
// __block_26
  end
  4'h4: begin
// __block_27_case
// __block_28
_d_readData = _w_p1hz_counter1hz;
// __block_29
  end
endcase
// __block_14
// __block_30
  end
  4'hf: begin
// __block_31_case
// __block_32
  case (in_memoryAddress[4+:4])
  4'h0: begin
// __block_34_case
// __block_35
  case (in_memoryAddress[0+:4])
  4'h7: begin
// __block_37_case
// __block_38
_d_readData = _w_gpu_processor_gpu_active;
// __block_39
  end
  4'h8: begin
// __block_40_case
// __block_41
_d_readData = _w_bitmap_window_bitmap_colour_read;
// __block_42
  end
endcase
// __block_36
// __block_43
  end
  4'h1: begin
// __block_44_case
// __block_45
  case (in_memoryAddress[0+:4])
  4'h5: begin
// __block_47_case
// __block_48
_d_readData = _w_character_map_window_tpu_active;
// __block_49
  end
endcase
// __block_46
// __block_50
  end
  4'h2: begin
// __block_51_case
// __block_52
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_54_case
// __block_55
_d_readData = _w_terminal_window_terminal_active;
// __block_56
  end
endcase
// __block_53
// __block_57
  end
  4'h3: begin
// __block_58_case
// __block_59
  case (in_memoryAddress[0+:4])
  4'h1: begin
// __block_61_case
// __block_62
_d_readData = _w_lower_sprites_sprite_read_active;
// __block_63
  end
  4'h2: begin
// __block_64_case
// __block_65
_d_readData = _w_lower_sprites_sprite_read_tile;
// __block_66
  end
  4'h3: begin
// __block_67_case
// __block_68
_d_readData = _w_lower_sprites_sprite_read_colour;
// __block_69
  end
  4'h4: begin
// __block_70_case
// __block_71
_d_readData = _w_lower_sprites_sprite_read_x;
// __block_72
  end
  4'h5: begin
// __block_73_case
// __block_74
_d_readData = _w_lower_sprites_sprite_read_y;
// __block_75
  end
  4'h6: begin
// __block_76_case
// __block_77
_d_readData = _w_lower_sprites_sprite_read_double;
// __block_78
  end
endcase
// __block_60
// __block_79
  end
  4'h4: begin
// __block_80_case
// __block_81
  case (in_memoryAddress[0+:4])
  4'h1: begin
// __block_83_case
// __block_84
_d_readData = _w_upper_sprites_sprite_read_active;
// __block_85
  end
  4'h2: begin
// __block_86_case
// __block_87
_d_readData = _w_upper_sprites_sprite_read_tile;
// __block_88
  end
  4'h3: begin
// __block_89_case
// __block_90
_d_readData = _w_upper_sprites_sprite_read_colour;
// __block_91
  end
  4'h4: begin
// __block_92_case
// __block_93
_d_readData = _w_upper_sprites_sprite_read_x;
// __block_94
  end
  4'h5: begin
// __block_95_case
// __block_96
_d_readData = _w_upper_sprites_sprite_read_y;
// __block_97
  end
  4'h6: begin
// __block_98_case
// __block_99
_d_readData = _w_upper_sprites_sprite_read_double;
// __block_100
  end
endcase
// __block_82
// __block_101
  end
  4'h5: begin
// __block_102_case
// __block_103
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_105_case
// __block_106
_d_readData = _w_lower_sprites_collision_0;
// __block_107
  end
  4'h1: begin
// __block_108_case
// __block_109
_d_readData = _w_lower_sprites_collision_1;
// __block_110
  end
  4'h2: begin
// __block_111_case
// __block_112
_d_readData = _w_lower_sprites_collision_2;
// __block_113
  end
  4'h3: begin
// __block_114_case
// __block_115
_d_readData = _w_lower_sprites_collision_3;
// __block_116
  end
  4'h4: begin
// __block_117_case
// __block_118
_d_readData = _w_lower_sprites_collision_4;
// __block_119
  end
  4'h5: begin
// __block_120_case
// __block_121
_d_readData = _w_lower_sprites_collision_5;
// __block_122
  end
  4'h6: begin
// __block_123_case
// __block_124
_d_readData = _w_lower_sprites_collision_6;
// __block_125
  end
  4'h7: begin
// __block_126_case
// __block_127
_d_readData = _w_lower_sprites_collision_7;
// __block_128
  end
  4'h8: begin
// __block_129_case
// __block_130
_d_readData = _w_lower_sprites_collision_8;
// __block_131
  end
  4'h9: begin
// __block_132_case
// __block_133
_d_readData = _w_lower_sprites_collision_9;
// __block_134
  end
  4'ha: begin
// __block_135_case
// __block_136
_d_readData = _w_lower_sprites_collision_10;
// __block_137
  end
  4'hb: begin
// __block_138_case
// __block_139
_d_readData = _w_lower_sprites_collision_11;
// __block_140
  end
  4'hc: begin
// __block_141_case
// __block_142
_d_readData = _w_lower_sprites_collision_12;
// __block_143
  end
endcase
// __block_104
// __block_144
  end
  4'h6: begin
// __block_145_case
// __block_146
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_148_case
// __block_149
_d_readData = _w_upper_sprites_collision_0;
// __block_150
  end
  4'h1: begin
// __block_151_case
// __block_152
_d_readData = _w_upper_sprites_collision_1;
// __block_153
  end
  4'h2: begin
// __block_154_case
// __block_155
_d_readData = _w_upper_sprites_collision_2;
// __block_156
  end
  4'h3: begin
// __block_157_case
// __block_158
_d_readData = _w_upper_sprites_collision_3;
// __block_159
  end
  4'h4: begin
// __block_160_case
// __block_161
_d_readData = _w_upper_sprites_collision_4;
// __block_162
  end
  4'h5: begin
// __block_163_case
// __block_164
_d_readData = _w_upper_sprites_collision_5;
// __block_165
  end
  4'h6: begin
// __block_166_case
// __block_167
_d_readData = _w_upper_sprites_collision_6;
// __block_168
  end
  4'h7: begin
// __block_169_case
// __block_170
_d_readData = _w_upper_sprites_collision_7;
// __block_171
  end
  4'h8: begin
// __block_172_case
// __block_173
_d_readData = _w_upper_sprites_collision_8;
// __block_174
  end
  4'h9: begin
// __block_175_case
// __block_176
_d_readData = _w_upper_sprites_collision_9;
// __block_177
  end
  4'ha: begin
// __block_178_case
// __block_179
_d_readData = _w_upper_sprites_collision_10;
// __block_180
  end
  4'hb: begin
// __block_181_case
// __block_182
_d_readData = _w_upper_sprites_collision_11;
// __block_183
  end
  4'hc: begin
// __block_184_case
// __block_185
_d_readData = _w_upper_sprites_collision_12;
// __block_186
  end
endcase
// __block_147
// __block_187
  end
  4'h7: begin
// __block_188_case
// __block_189
  case (in_memoryAddress[0+:4])
  4'h4: begin
// __block_191_case
// __block_192
_d_readData = _w_gpu_processor_vector_block_active;
// __block_193
  end
endcase
// __block_190
// __block_194
  end
  4'h9: begin
// __block_195_case
// __block_196
  case (in_memoryAddress[0+:4])
  4'h9: begin
// __block_198_case
// __block_199
_d_readData = _w_tile_map_tm_lastaction;
// __block_200
  end
  4'ha: begin
// __block_201_case
// __block_202
_d_readData = _w_tile_map_tm_active;
// __block_203
  end
endcase
// __block_197
// __block_204
  end
  4'ha: begin
// __block_205_case
// __block_206
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_208_case
// __block_209
_d_readData = _w_doperations2_total[16+:16];
// __block_210
  end
  4'h1: begin
// __block_211_case
// __block_212
_d_readData = _w_doperations2_total[0+:16];
// __block_213
  end
  4'h2: begin
// __block_214_case
// __block_215
_d_readData = _w_doperations2_difference[16+:16];
// __block_216
  end
  4'h3: begin
// __block_217_case
// __block_218
_d_readData = _w_doperations2_difference[0+:16];
// __block_219
  end
  4'h4: begin
// __block_220_case
// __block_221
_d_readData = _w_doperations1_increment[16+:16];
// __block_222
  end
  4'h5: begin
// __block_223_case
// __block_224
_d_readData = _w_doperations1_increment[0+:16];
// __block_225
  end
  4'h6: begin
// __block_226_case
// __block_227
_d_readData = _w_doperations1_decrement[16+:16];
// __block_228
  end
  4'h7: begin
// __block_229_case
// __block_230
_d_readData = _w_doperations1_decrement[0+:16];
// __block_231
  end
  4'h8: begin
// __block_232_case
// __block_233
_d_readData = _w_doperations1_times2[16+:16];
// __block_234
  end
  4'h9: begin
// __block_235_case
// __block_236
_d_readData = _w_doperations1_times2[0+:16];
// __block_237
  end
  4'ha: begin
// __block_238_case
// __block_239
_d_readData = _w_doperations1_divide2[16+:16];
// __block_240
  end
  4'hb: begin
// __block_241_case
// __block_242
_d_readData = _w_doperations1_divide2[0+:16];
// __block_243
  end
  4'hc: begin
// __block_244_case
// __block_245
_d_readData = _w_doperations1_negation[16+:16];
// __block_246
  end
  4'hd: begin
// __block_247_case
// __block_248
_d_readData = _w_doperations1_negation[0+:16];
// __block_249
  end
  4'he: begin
// __block_250_case
// __block_251
_d_readData = _w_doperations1_binaryinvert[16+:16];
// __block_252
  end
  4'hf: begin
// __block_253_case
// __block_254
_d_readData = _w_doperations1_binaryinvert[0+:16];
// __block_255
  end
endcase
// __block_207
// __block_256
  end
  4'hb: begin
// __block_257_case
// __block_258
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_260_case
// __block_261
_d_readData = _w_doperations2_binaryxor[16+:16];
// __block_262
  end
  4'h1: begin
// __block_263_case
// __block_264
_d_readData = _w_doperations2_binaryxor[0+:16];
// __block_265
  end
  4'h2: begin
// __block_266_case
// __block_267
_d_readData = _w_doperations2_binaryand[16+:16];
// __block_268
  end
  4'h3: begin
// __block_269_case
// __block_270
_d_readData = _w_doperations2_binaryand[0+:16];
// __block_271
  end
  4'h4: begin
// __block_272_case
// __block_273
_d_readData = _w_doperations2_binaryor[16+:16];
// __block_274
  end
  4'h5: begin
// __block_275_case
// __block_276
_d_readData = _w_doperations2_binaryor[0+:16];
// __block_277
  end
  4'h6: begin
// __block_278_case
// __block_279
_d_readData = _w_doperations1_absolute[16+:16];
// __block_280
  end
  4'h7: begin
// __block_281_case
// __block_282
_d_readData = _w_doperations1_absolute[0+:16];
// __block_283
  end
  4'h8: begin
// __block_284_case
// __block_285
_d_readData = _w_doperations2_maximum[16+:16];
// __block_286
  end
  4'h9: begin
// __block_287_case
// __block_288
_d_readData = _w_doperations2_maximum[0+:16];
// __block_289
  end
  4'ha: begin
// __block_290_case
// __block_291
_d_readData = _w_doperations2_minimum[16+:16];
// __block_292
  end
  4'hb: begin
// __block_293_case
// __block_294
_d_readData = _w_doperations2_minimum[0+:16];
// __block_295
  end
  4'hc: begin
// __block_296_case
// __block_297
_d_readData = _w_doperations1_zeroequal;
// __block_298
  end
  4'hd: begin
// __block_299_case
// __block_300
_d_readData = _w_doperations1_zeroless;
// __block_301
  end
  4'he: begin
// __block_302_case
// __block_303
_d_readData = _w_doperations2_equal;
// __block_304
  end
  4'hf: begin
// __block_305_case
// __block_306
_d_readData = _w_doperations2_lessthan;
// __block_307
  end
endcase
// __block_259
// __block_308
  end
  4'hd: begin
// __block_309_case
// __block_310
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_312_case
// __block_313
_d_readData = _w_divmod32by16to16qr_quotient[0+:16];
// __block_314
  end
  4'h1: begin
// __block_315_case
// __block_316
_d_readData = _w_divmod32by16to16qr_remainder[0+:16];
// __block_317
  end
  4'h3: begin
// __block_318_case
// __block_319
_d_readData = _w_divmod32by16to16qr_active;
// __block_320
  end
  4'h4: begin
// __block_321_case
// __block_322
_d_readData = _w_divmod16by16to16qr_quotient;
// __block_323
  end
  4'h5: begin
// __block_324_case
// __block_325
_d_readData = _w_divmod16by16to16qr_remainder;
// __block_326
  end
  4'h6: begin
// __block_327_case
// __block_328
_d_readData = _w_divmod16by16to16qr_active;
// __block_329
  end
  4'h7: begin
// __block_330_case
// __block_331
_d_readData = _w_multiplier16by16to32_product[16+:16];
// __block_332
  end
  4'h8: begin
// __block_333_case
// __block_334
_d_readData = _w_multiplier16by16to32_product[0+:16];
// __block_335
  end
  4'h9: begin
// __block_336_case
// __block_337
_d_readData = _w_multiplier16by16to32_active;
// __block_338
  end
endcase
// __block_311
// __block_339
  end
  4'he: begin
// __block_340_case
// __block_341
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_343_case
// __block_344
_d_readData = _w_rng_g_noise_out;
// __block_345
  end
  4'h3: begin
// __block_346_case
// __block_347
_d_readData = _w_apu_processor_L_audio_active;
// __block_348
  end
  4'h7: begin
// __block_349_case
// __block_350
_d_readData = _w_apu_processor_R_audio_active;
// __block_351
  end
  4'hd: begin
// __block_352_case
// __block_353
_d_readData = _w_timer1hz_counter1hz;
// __block_354
  end
  4'he: begin
// __block_355_case
// __block_356
_d_readData = _w_timer1khz_counter1khz;
// __block_357
  end
  4'hf: begin
// __block_358_case
// __block_359
_d_readData = _w_sleepTimer_counter1khz;
// __block_360
  end
endcase
// __block_342
// __block_361
  end
  4'hf: begin
// __block_362_case
// __block_363
  case (in_memoryAddress[0+:4])
  4'hf: begin
// __block_365_case
// __block_366
_d_readData = in_vblank;
// __block_367
  end
endcase
// __block_364
// __block_368
  end
endcase
// __block_33
// __block_369
  end
endcase
// __block_11
// __block_370
  end
endcase
// __block_8
// __block_371
end else begin
// __block_6
end
// __block_372
if (in_memoryWrite) begin
// __block_373
// __block_375
_d_coProReset = 3;
  case (in_memoryAddress[12+:4])
  4'hf: begin
// __block_377_case
// __block_378
  case (in_memoryAddress[8+:4])
  4'h0: begin
// __block_380_case
// __block_381
  case (in_memoryAddress[0+:4])
  4'h0: begin
// __block_383_case
// __block_384
_d_uartOutBuffer_wdata1 = in_writeData[0+:8];
_d_newuartOutBufferTop = _d_uartOutBufferTop+1;
// __block_385
  end
  4'h2: begin
// __block_386_case
// __block_387
_d_leds = in_writeData;
// __block_388
  end
endcase
// __block_382
// __block_389
  end
  4'hf: begin
// __block_390_case
// __block_391
  case (in_memoryAddress[0+:8])
  8'h00: begin
// __block_393_case
// __block_394
_d_gpu_processor_gpu_x = in_writeData;
// __block_395
  end
  8'h01: begin
// __block_396_case
// __block_397
_d_gpu_processor_gpu_y = in_writeData;
// __block_398
  end
  8'h02: begin
// __block_399_case
// __block_400
_d_gpu_processor_gpu_colour = in_writeData;
// __block_401
  end
  8'h03: begin
// __block_402_case
// __block_403
_d_gpu_processor_gpu_param0 = in_writeData;
// __block_404
  end
  8'h04: begin
// __block_405_case
// __block_406
_d_gpu_processor_gpu_param1 = in_writeData;
// __block_407
  end
  8'h05: begin
// __block_408_case
// __block_409
_d_gpu_processor_gpu_param2 = in_writeData;
// __block_410
  end
  8'h06: begin
// __block_411_case
// __block_412
_d_gpu_processor_gpu_param3 = in_writeData;
// __block_413
  end
  8'h07: begin
// __block_414_case
// __block_415
_d_gpu_processor_gpu_write = in_writeData;
// __block_416
  end
  8'h08: begin
// __block_417_case
// __block_418
_d_bitmap_window_bitmap_write_offset = in_writeData;
// __block_419
  end
  8'h09: begin
// __block_420_case
// __block_421
_d_bitmap_window_bitmap_x_read = in_writeData;
// __block_422
  end
  8'h0a: begin
// __block_423_case
// __block_424
_d_bitmap_window_bitmap_y_read = in_writeData;
// __block_425
  end
  8'h0b: begin
// __block_426_case
// __block_427
_d_gpu_processor_blit1_writer_tile = in_writeData;
// __block_428
  end
  8'h0c: begin
// __block_429_case
// __block_430
_d_gpu_processor_blit1_writer_line = in_writeData;
// __block_431
  end
  8'h0d: begin
// __block_432_case
// __block_433
_d_gpu_processor_blit1_writer_bitmap = in_writeData;
// __block_434
  end
  8'h10: begin
// __block_435_case
// __block_436
_d_character_map_window_tpu_x = in_writeData;
// __block_437
  end
  8'h11: begin
// __block_438_case
// __block_439
_d_character_map_window_tpu_y = in_writeData;
// __block_440
  end
  8'h12: begin
// __block_441_case
// __block_442
_d_character_map_window_tpu_character = in_writeData;
// __block_443
  end
  8'h13: begin
// __block_444_case
// __block_445
_d_character_map_window_tpu_background = in_writeData;
// __block_446
  end
  8'h14: begin
// __block_447_case
// __block_448
_d_character_map_window_tpu_foreground = in_writeData;
// __block_449
  end
  8'h15: begin
// __block_450_case
// __block_451
_d_character_map_window_tpu_write = in_writeData;
// __block_452
  end
  8'h20: begin
// __block_453_case
// __block_454
_d_terminal_window_terminal_character = in_writeData;
_d_terminal_window_terminal_write = 1;
// __block_455
  end
  8'h21: begin
// __block_456_case
// __block_457
_d_terminal_window_showterminal = in_writeData;
// __block_458
  end
  8'h30: begin
// __block_459_case
// __block_460
_d_lower_sprites_sprite_set_number = in_writeData;
// __block_461
  end
  8'h31: begin
// __block_462_case
// __block_463
_d_lower_sprites_sprite_set_active = in_writeData;
_d_lower_sprites_sprite_layer_write = 1;
// __block_464
  end
  8'h32: begin
// __block_465_case
// __block_466
_d_lower_sprites_sprite_set_tile = in_writeData;
_d_lower_sprites_sprite_layer_write = 2;
// __block_467
  end
  8'h33: begin
// __block_468_case
// __block_469
_d_lower_sprites_sprite_set_colour = in_writeData;
_d_lower_sprites_sprite_layer_write = 3;
// __block_470
  end
  8'h34: begin
// __block_471_case
// __block_472
_d_lower_sprites_sprite_set_x = in_writeData;
_d_lower_sprites_sprite_layer_write = 4;
// __block_473
  end
  8'h35: begin
// __block_474_case
// __block_475
_d_lower_sprites_sprite_set_y = in_writeData;
_d_lower_sprites_sprite_layer_write = 5;
// __block_476
  end
  8'h36: begin
// __block_477_case
// __block_478
_d_lower_sprites_sprite_set_double = in_writeData;
_d_lower_sprites_sprite_layer_write = 6;
// __block_479
  end
  8'h38: begin
// __block_480_case
// __block_481
_d_lower_sprites_sprite_writer_sprite = in_writeData;
// __block_482
  end
  8'h39: begin
// __block_483_case
// __block_484
_d_lower_sprites_sprite_writer_line = in_writeData;
// __block_485
  end
  8'h3a: begin
// __block_486_case
// __block_487
_d_lower_sprites_sprite_writer_bitmap = in_writeData;
_d_lower_sprites_sprite_writer_active = 1;
// __block_488
  end
  8'h3e: begin
// __block_489_case
// __block_490
_d_lower_sprites_sprite_update = in_writeData;
_d_lower_sprites_sprite_layer_write = 10;
// __block_491
  end
  8'h40: begin
// __block_492_case
// __block_493
_d_upper_sprites_sprite_set_number = in_writeData;
// __block_494
  end
  8'h41: begin
// __block_495_case
// __block_496
_d_upper_sprites_sprite_set_active = in_writeData;
_d_upper_sprites_sprite_layer_write = 1;
// __block_497
  end
  8'h42: begin
// __block_498_case
// __block_499
_d_upper_sprites_sprite_set_tile = in_writeData;
_d_upper_sprites_sprite_layer_write = 2;
// __block_500
  end
  8'h43: begin
// __block_501_case
// __block_502
_d_upper_sprites_sprite_set_colour = in_writeData;
_d_upper_sprites_sprite_layer_write = 3;
// __block_503
  end
  8'h44: begin
// __block_504_case
// __block_505
_d_upper_sprites_sprite_set_x = in_writeData;
_d_upper_sprites_sprite_layer_write = 4;
// __block_506
  end
  8'h45: begin
// __block_507_case
// __block_508
_d_upper_sprites_sprite_set_y = in_writeData;
_d_upper_sprites_sprite_layer_write = 5;
// __block_509
  end
  8'h46: begin
// __block_510_case
// __block_511
_d_upper_sprites_sprite_set_double = in_writeData;
_d_upper_sprites_sprite_layer_write = 6;
// __block_512
  end
  8'h48: begin
// __block_513_case
// __block_514
_d_upper_sprites_sprite_writer_sprite = in_writeData;
// __block_515
  end
  8'h49: begin
// __block_516_case
// __block_517
_d_upper_sprites_sprite_writer_line = in_writeData;
// __block_518
  end
  8'h4a: begin
// __block_519_case
// __block_520
_d_upper_sprites_sprite_writer_bitmap = in_writeData;
_d_upper_sprites_sprite_writer_active = 1;
// __block_521
  end
  8'h4e: begin
// __block_522_case
// __block_523
_d_upper_sprites_sprite_update = in_writeData;
_d_upper_sprites_sprite_layer_write = 10;
// __block_524
  end
  8'h70: begin
// __block_525_case
// __block_526
_d_gpu_processor_vector_block_number = in_writeData;
// __block_527
  end
  8'h71: begin
// __block_528_case
// __block_529
_d_gpu_processor_vector_block_colour = in_writeData;
// __block_530
  end
  8'h72: begin
// __block_531_case
// __block_532
_d_gpu_processor_vector_block_xc = in_writeData;
// __block_533
  end
  8'h73: begin
// __block_534_case
// __block_535
_d_gpu_processor_vector_block_yc = in_writeData;
// __block_536
  end
  8'h74: begin
// __block_537_case
// __block_538
_d_gpu_processor_draw_vector = 1;
// __block_539
  end
  8'h75: begin
// __block_540_case
// __block_541
_d_gpu_processor_vertices_writer_block = in_writeData;
// __block_542
  end
  8'h76: begin
// __block_543_case
// __block_544
_d_gpu_processor_vertices_writer_vertex = in_writeData;
// __block_545
  end
  8'h77: begin
// __block_546_case
// __block_547
_d_gpu_processor_vertices_writer_xdelta = in_writeData;
// __block_548
  end
  8'h78: begin
// __block_549_case
// __block_550
_d_gpu_processor_vertices_writer_ydelta = in_writeData;
// __block_551
  end
  8'h79: begin
// __block_552_case
// __block_553
_d_gpu_processor_vertices_writer_active = in_writeData;
// __block_554
  end
  8'h90: begin
// __block_555_case
// __block_556
_d_tile_map_tm_x = in_writeData;
// __block_557
  end
  8'h91: begin
// __block_558_case
// __block_559
_d_tile_map_tm_y = in_writeData;
// __block_560
  end
  8'h92: begin
// __block_561_case
// __block_562
_d_tile_map_tm_character = in_writeData;
// __block_563
  end
  8'h93: begin
// __block_564_case
// __block_565
_d_tile_map_tm_background = in_writeData;
// __block_566
  end
  8'h94: begin
// __block_567_case
// __block_568
_d_tile_map_tm_foreground = in_writeData;
// __block_569
  end
  8'h95: begin
// __block_570_case
// __block_571
_d_tile_map_tm_write = 1;
// __block_572
  end
  8'h96: begin
// __block_573_case
// __block_574
_d_tile_map_tile_writer_tile = in_writeData;
// __block_575
  end
  8'h97: begin
// __block_576_case
// __block_577
_d_tile_map_tile_writer_line = in_writeData;
// __block_578
  end
  8'h98: begin
// __block_579_case
// __block_580
_d_tile_map_tile_writer_bitmap = in_writeData;
// __block_581
  end
  8'h99: begin
// __block_582_case
// __block_583
_d_tile_map_tm_scrollwrap = in_writeData;
// __block_584
  end
  8'ha0: begin
// __block_585_case
// __block_586
_d_doperations2_operand1h = in_writeData;
_d_doperations1_operand1h = in_writeData;
// __block_587
  end
  8'ha1: begin
// __block_588_case
// __block_589
_d_doperations2_operand1l = in_writeData;
_d_doperations1_operand1l = in_writeData;
// __block_590
  end
  8'ha2: begin
// __block_591_case
// __block_592
_d_doperations2_operand2h = in_writeData;
// __block_593
  end
  8'ha3: begin
// __block_594_case
// __block_595
_d_doperations2_operand2l = in_writeData;
// __block_596
  end
  8'hd0: begin
// __block_597_case
// __block_598
_d_divmod32by16to16qr_dividendh = in_writeData;
// __block_599
  end
  8'hd1: begin
// __block_600_case
// __block_601
_d_divmod32by16to16qr_dividendl = in_writeData;
// __block_602
  end
  8'hd2: begin
// __block_603_case
// __block_604
_d_divmod32by16to16qr_divisor = in_writeData;
// __block_605
  end
  8'hd3: begin
// __block_606_case
// __block_607
_d_divmod32by16to16qr_start = in_writeData;
// __block_608
  end
  8'hd4: begin
// __block_609_case
// __block_610
_d_divmod16by16to16qr_dividend = in_writeData;
// __block_611
  end
  8'hd5: begin
// __block_612_case
// __block_613
_d_divmod16by16to16qr_divisor = in_writeData;
// __block_614
  end
  8'hd6: begin
// __block_615_case
// __block_616
_d_divmod16by16to16qr_start = in_writeData;
// __block_617
  end
  8'hd7: begin
// __block_618_case
// __block_619
_d_multiplier16by16to32_factor1 = in_writeData;
// __block_620
  end
  8'hd8: begin
// __block_621_case
// __block_622
_d_multiplier16by16to32_factor2 = in_writeData;
// __block_623
  end
  8'hd9: begin
// __block_624_case
// __block_625
_d_multiplier16by16to32_start = in_writeData;
// __block_626
  end
  8'he0: begin
// __block_627_case
// __block_628
_d_apu_processor_L_waveform = in_writeData;
// __block_629
  end
  8'he1: begin
// __block_630_case
// __block_631
_d_apu_processor_L_note = in_writeData;
// __block_632
  end
  8'he2: begin
// __block_633_case
// __block_634
_d_apu_processor_L_duration = in_writeData;
// __block_635
  end
  8'he3: begin
// __block_636_case
// __block_637
_d_apu_processor_L_apu_write = in_writeData;
// __block_638
  end
  8'he4: begin
// __block_639_case
// __block_640
_d_apu_processor_R_waveform = in_writeData;
// __block_641
  end
  8'he5: begin
// __block_642_case
// __block_643
_d_apu_processor_R_note = in_writeData;
// __block_644
  end
  8'he6: begin
// __block_645_case
// __block_646
_d_apu_processor_R_duration = in_writeData;
// __block_647
  end
  8'he7: begin
// __block_648_case
// __block_649
_d_apu_processor_R_apu_write = in_writeData;
// __block_650
  end
  8'he8: begin
// __block_651_case
// __block_652
_d_rng_resetRandom = 1;
// __block_653
  end
  8'hed: begin
// __block_654_case
// __block_655
_d_timer1hz_resetCounter = 1;
// __block_656
  end
  8'hee: begin
// __block_657_case
// __block_658
_d_timer1khz_resetCount = in_writeData;
_d_timer1khz_resetCounter = 1;
// __block_659
  end
  8'hef: begin
// __block_660_case
// __block_661
_d_sleepTimer_resetCount = in_writeData;
_d_sleepTimer_resetCounter = 1;
// __block_662
  end
  8'hf0: begin
// __block_663_case
// __block_664
_d_background_generator_backgroundcolour = in_writeData;
_d_background_generator_background_write = 1;
// __block_665
  end
  8'hf1: begin
// __block_666_case
// __block_667
_d_background_generator_backgroundcolour_alt = in_writeData;
_d_background_generator_background_write = 2;
// __block_668
  end
  8'hf2: begin
// __block_669_case
// __block_670
_d_background_generator_backgroundcolour_mode = in_writeData;
_d_background_generator_background_write = 3;
// __block_671
  end
endcase
// __block_392
// __block_672
  end
endcase
// __block_379
// __block_673
  end
endcase
// __block_376
// __block_674
end else begin
// __block_374
// __block_675
_d_coProReset = (_q_coProReset==0)?0:_q_coProReset-1;
// __block_676
end
// __block_677
if (_d_coProReset==1) begin
// __block_678
// __block_680
_d_background_generator_background_write = 0;
_d_tile_map_tm_write = 0;
_d_tile_map_tm_scrollwrap = 0;
_d_lower_sprites_sprite_layer_write = 0;
_d_lower_sprites_sprite_writer_active = 0;
_d_bitmap_window_bitmap_write_offset = 0;
_d_gpu_processor_gpu_write = 0;
_d_gpu_processor_draw_vector = 0;
_d_upper_sprites_sprite_layer_write = 0;
_d_upper_sprites_sprite_writer_active = 0;
_d_character_map_window_tpu_write = 0;
_d_terminal_window_terminal_write = 0;
_d_apu_processor_L_apu_write = 0;
_d_apu_processor_R_apu_write = 0;
// __block_681
end else begin
// __block_679
end
// __block_682
// __block_683
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of memmap_io
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_main_mem_dstack(
input      [7:0]                in_dstack_addr0,
output reg  [15:0]     out_dstack_rdata0,
output reg  [15:0]     out_dstack_rdata1,
input      [0:0]             in_dstack_wenable1,
input      [15:0]                 in_dstack_wdata1,
input      [7:0]                in_dstack_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[255:0];
always @(posedge clock0) begin
  out_dstack_rdata0 <= buffer[in_dstack_addr0];
end
always @(posedge clock1) begin
  if (in_dstack_wenable1) begin
    buffer[in_dstack_addr1] <= in_dstack_wdata1;
  end
end

endmodule

module M_main_mem_rstack(
input      [7:0]                in_rstack_addr0,
output reg  [15:0]     out_rstack_rdata0,
output reg  [15:0]     out_rstack_rdata1,
input      [0:0]             in_rstack_wenable1,
input      [15:0]                 in_rstack_wdata1,
input      [7:0]                in_rstack_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[255:0];
always @(posedge clock0) begin
  out_rstack_rdata0 <= buffer[in_rstack_addr0];
end
always @(posedge clock1) begin
  if (in_rstack_wenable1) begin
    buffer[in_rstack_addr1] <= in_rstack_wdata1;
  end
end

endmodule

module M_main_mem_ram(
input      [13:0]                in_ram_addr0,
output reg  [15:0]     out_ram_rdata0,
output reg  [15:0]     out_ram_rdata1,
input      [0:0]             in_ram_wenable1,
input      [15:0]                 in_ram_wdata1,
input      [13:0]                in_ram_addr1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[16383:0];
always @(posedge clock0) begin
  out_ram_rdata0 <= buffer[in_ram_addr0];
end
always @(posedge clock1) begin
  if (in_ram_wenable1) begin
    buffer[in_ram_addr1] <= in_ram_wdata1;
  end
end
initial begin
 buffer[0] = 16'h0CF0;
 buffer[1] = 16'h0010;
 buffer[2] = 16'h0000;
 buffer[3] = 16'h0000;
 buffer[4] = 16'h0000;
 buffer[5] = 16'h7F00;
 buffer[6] = 16'h0E24;
 buffer[7] = 16'h0F02;
 buffer[8] = 16'h0000;
 buffer[9] = 16'h0000;
 buffer[10] = 16'h0000;
 buffer[11] = 16'h0000;
 buffer[12] = 16'h0000;
 buffer[13] = 16'h0000;
 buffer[14] = 16'h0000;
 buffer[15] = 16'h0000;
 buffer[16] = 16'h2406;
 buffer[17] = 16'h23EE;
 buffer[18] = 16'h0940;
 buffer[19] = 16'h0952;
 buffer[20] = 16'h19A8;
 buffer[21] = 16'h0BE0;
 buffer[22] = 16'h0CCC;
 buffer[23] = 16'h13D8;
 buffer[24] = 16'h145A;
 buffer[25] = 16'h1482;
 buffer[26] = 16'h14EE;
 buffer[27] = 16'h0000;
 buffer[28] = 16'h0000;
 buffer[29] = 16'h0000;
 buffer[30] = 16'h0000;
 buffer[31] = 16'h0000;
 buffer[32] = 16'h0000;
 buffer[33] = 16'h0000;
 buffer[34] = 16'h0000;
 buffer[35] = 16'h0000;
 buffer[36] = 16'h0000;
 buffer[37] = 16'h0000;
 buffer[38] = 16'h0000;
 buffer[39] = 16'h0000;
 buffer[40] = 16'h0000;
 buffer[41] = 16'h0000;
 buffer[42] = 16'h0000;
 buffer[43] = 16'h0000;
 buffer[44] = 16'h0000;
 buffer[45] = 16'h0000;
 buffer[46] = 16'h0000;
 buffer[47] = 16'h0000;
 buffer[48] = 16'h0000;
 buffer[49] = 16'h0000;
 buffer[50] = 16'h0000;
 buffer[51] = 16'h0000;
 buffer[52] = 16'h0000;
 buffer[53] = 16'h0000;
 buffer[54] = 16'h0000;
 buffer[55] = 16'h0000;
 buffer[56] = 16'h0000;
 buffer[57] = 16'h0000;
 buffer[58] = 16'h0000;
 buffer[59] = 16'h0000;
 buffer[60] = 16'h0000;
 buffer[61] = 16'h0000;
 buffer[62] = 16'h0000;
 buffer[63] = 16'h0000;
 buffer[64] = 16'h6003;
 buffer[65] = 16'h6003;
 buffer[66] = 16'h6003;
 buffer[67] = 16'h6003;
 buffer[68] = 16'h6003;
 buffer[69] = 16'h6003;
 buffer[70] = 16'h6003;
 buffer[71] = 16'h6003;
 buffer[72] = 16'h6003;
 buffer[73] = 16'h6003;
 buffer[74] = 16'h6003;
 buffer[75] = 16'h6003;
 buffer[76] = 16'h6003;
 buffer[77] = 16'h6003;
 buffer[78] = 16'h6003;
 buffer[79] = 16'h710C;
 buffer[80] = 16'h6001;
 buffer[81] = 16'h6001;
 buffer[82] = 16'h6001;
 buffer[83] = 16'h6001;
 buffer[84] = 16'h6001;
 buffer[85] = 16'h6001;
 buffer[86] = 16'h6001;
 buffer[87] = 16'h6001;
 buffer[88] = 16'h6001;
 buffer[89] = 16'h6001;
 buffer[90] = 16'h6001;
 buffer[91] = 16'h6001;
 buffer[92] = 16'h6001;
 buffer[93] = 16'h6001;
 buffer[94] = 16'h6001;
 buffer[95] = 16'h700C;
 buffer[96] = 16'h6100;
 buffer[97] = 16'h700C;
 buffer[98] = 16'h404E;
 buffer[99] = 16'h005E;
 buffer[100] = 16'h404D;
 buffer[101] = 16'h005D;
 buffer[102] = 16'h404C;
 buffer[103] = 16'h005C;
 buffer[104] = 16'h404B;
 buffer[105] = 16'h005B;
 buffer[106] = 16'h404A;
 buffer[107] = 16'h005A;
 buffer[108] = 16'h4049;
 buffer[109] = 16'h0059;
 buffer[110] = 16'h4048;
 buffer[111] = 16'h0058;
 buffer[112] = 16'h4047;
 buffer[113] = 16'h0057;
 buffer[114] = 16'h4046;
 buffer[115] = 16'h0056;
 buffer[116] = 16'h4045;
 buffer[117] = 16'h0055;
 buffer[118] = 16'h4044;
 buffer[119] = 16'h0054;
 buffer[120] = 16'h4043;
 buffer[121] = 16'h0053;
 buffer[122] = 16'h4042;
 buffer[123] = 16'h0052;
 buffer[124] = 16'h4041;
 buffer[125] = 16'h0051;
 buffer[126] = 16'h4040;
 buffer[127] = 16'h0050;
 buffer[128] = 16'h700C;
 buffer[129] = 16'h0000;
 buffer[130] = 16'h0000;
 buffer[131] = 16'h0000;
 buffer[132] = 16'h0000;
 buffer[133] = 16'h0000;
 buffer[134] = 16'h0000;
 buffer[135] = 16'h0000;
 buffer[136] = 16'h0000;
 buffer[137] = 16'h0000;
 buffer[138] = 16'h0000;
 buffer[139] = 16'h0000;
 buffer[140] = 16'h0000;
 buffer[141] = 16'h0000;
 buffer[142] = 16'h0000;
 buffer[143] = 16'h0000;
 buffer[144] = 16'h0000;
 buffer[145] = 16'h0000;
 buffer[146] = 16'h0000;
 buffer[147] = 16'h0000;
 buffer[148] = 16'h0000;
 buffer[149] = 16'h0000;
 buffer[150] = 16'h0000;
 buffer[151] = 16'h0000;
 buffer[152] = 16'h0000;
 buffer[153] = 16'h0000;
 buffer[154] = 16'h0000;
 buffer[155] = 16'h0000;
 buffer[156] = 16'h0000;
 buffer[157] = 16'h0000;
 buffer[158] = 16'h0000;
 buffer[159] = 16'h0000;
 buffer[160] = 16'h0000;
 buffer[161] = 16'h0000;
 buffer[162] = 16'h0000;
 buffer[163] = 16'h0000;
 buffer[164] = 16'h0000;
 buffer[165] = 16'h0000;
 buffer[166] = 16'h0000;
 buffer[167] = 16'h0000;
 buffer[168] = 16'h0000;
 buffer[169] = 16'h0000;
 buffer[170] = 16'h0000;
 buffer[171] = 16'h0000;
 buffer[172] = 16'h0000;
 buffer[173] = 16'h0000;
 buffer[174] = 16'h0000;
 buffer[175] = 16'h0000;
 buffer[176] = 16'h0000;
 buffer[177] = 16'h0000;
 buffer[178] = 16'h0000;
 buffer[179] = 16'h0000;
 buffer[180] = 16'h0000;
 buffer[181] = 16'h0000;
 buffer[182] = 16'h0000;
 buffer[183] = 16'h0000;
 buffer[184] = 16'h0000;
 buffer[185] = 16'h0000;
 buffer[186] = 16'h0000;
 buffer[187] = 16'h0000;
 buffer[188] = 16'h0000;
 buffer[189] = 16'h0000;
 buffer[190] = 16'h0000;
 buffer[191] = 16'h0000;
 buffer[192] = 16'h0000;
 buffer[193] = 16'h6E04;
 buffer[194] = 16'h6F6F;
 buffer[195] = 16'h0070;
 buffer[196] = 16'h700C;
 buffer[197] = 16'h0182;
 buffer[198] = 16'h2B01;
 buffer[199] = 16'h720F;
 buffer[200] = 16'h018C;
 buffer[201] = 16'h7803;
 buffer[202] = 16'h726F;
 buffer[203] = 16'h750F;
 buffer[204] = 16'h0192;
 buffer[205] = 16'h6103;
 buffer[206] = 16'h646E;
 buffer[207] = 16'h730F;
 buffer[208] = 16'h019A;
 buffer[209] = 16'h6F02;
 buffer[210] = 16'h0072;
 buffer[211] = 16'h740F;
 buffer[212] = 16'h01A2;
 buffer[213] = 16'h6906;
 buffer[214] = 16'h766E;
 buffer[215] = 16'h7265;
 buffer[216] = 16'h0074;
 buffer[217] = 16'h760C;
 buffer[218] = 16'h01AA;
 buffer[219] = 16'h3D01;
 buffer[220] = 16'h770F;
 buffer[221] = 16'h01B6;
 buffer[222] = 16'h3C01;
 buffer[223] = 16'h780F;
 buffer[224] = 16'h01BC;
 buffer[225] = 16'h7502;
 buffer[226] = 16'h003C;
 buffer[227] = 16'h7F0F;
 buffer[228] = 16'h01C2;
 buffer[229] = 16'h7304;
 buffer[230] = 16'h6177;
 buffer[231] = 16'h0070;
 buffer[232] = 16'h718C;
 buffer[233] = 16'h01CA;
 buffer[234] = 16'h7502;
 buffer[235] = 16'h003E;
 buffer[236] = 16'h6180;
 buffer[237] = 16'h7F0F;
 buffer[238] = 16'h01D4;
 buffer[239] = 16'h6403;
 buffer[240] = 16'h7075;
 buffer[241] = 16'h708D;
 buffer[242] = 16'h01DE;
 buffer[243] = 16'h6404;
 buffer[244] = 16'h6F72;
 buffer[245] = 16'h0070;
 buffer[246] = 16'h710F;
 buffer[247] = 16'h01E6;
 buffer[248] = 16'h6F04;
 buffer[249] = 16'h6576;
 buffer[250] = 16'h0072;
 buffer[251] = 16'h718D;
 buffer[252] = 16'h01F0;
 buffer[253] = 16'h6E03;
 buffer[254] = 16'h7069;
 buffer[255] = 16'h700F;
 buffer[256] = 16'h01FA;
 buffer[257] = 16'h6C06;
 buffer[258] = 16'h6873;
 buffer[259] = 16'h6669;
 buffer[260] = 16'h0074;
 buffer[261] = 16'h7D0F;
 buffer[262] = 16'h0202;
 buffer[263] = 16'h7206;
 buffer[264] = 16'h6873;
 buffer[265] = 16'h6669;
 buffer[266] = 16'h0074;
 buffer[267] = 16'h790F;
 buffer[268] = 16'h020E;
 buffer[269] = 16'h3102;
 buffer[270] = 16'h002D;
 buffer[271] = 16'h7A0C;
 buffer[272] = 16'h021A;
 buffer[273] = 16'h3E42;
 buffer[274] = 16'h0072;
 buffer[275] = 16'h6B8D;
 buffer[276] = 16'h6180;
 buffer[277] = 16'h6147;
 buffer[278] = 16'h6147;
 buffer[279] = 16'h700C;
 buffer[280] = 16'h0222;
 buffer[281] = 16'h7242;
 buffer[282] = 16'h003E;
 buffer[283] = 16'h6B8D;
 buffer[284] = 16'h6B8D;
 buffer[285] = 16'h6180;
 buffer[286] = 16'h6147;
 buffer[287] = 16'h700C;
 buffer[288] = 16'h0232;
 buffer[289] = 16'h7242;
 buffer[290] = 16'h0040;
 buffer[291] = 16'h6B8D;
 buffer[292] = 16'h6B8D;
 buffer[293] = 16'h6081;
 buffer[294] = 16'h6147;
 buffer[295] = 16'h6180;
 buffer[296] = 16'h6147;
 buffer[297] = 16'h700C;
 buffer[298] = 16'h0242;
 buffer[299] = 16'h4001;
 buffer[300] = 16'h7C0C;
 buffer[301] = 16'h0256;
 buffer[302] = 16'h2101;
 buffer[303] = 16'h6023;
 buffer[304] = 16'h710F;
 buffer[305] = 16'h025C;
 buffer[306] = 16'h3C02;
 buffer[307] = 16'h003E;
 buffer[308] = 16'h721F;
 buffer[309] = 16'h0264;
 buffer[310] = 16'h3002;
 buffer[311] = 16'h003C;
 buffer[312] = 16'h791C;
 buffer[313] = 16'h026C;
 buffer[314] = 16'h3002;
 buffer[315] = 16'h003D;
 buffer[316] = 16'h701C;
 buffer[317] = 16'h0274;
 buffer[318] = 16'h3003;
 buffer[319] = 16'h3E3C;
 buffer[320] = 16'h711C;
 buffer[321] = 16'h027C;
 buffer[322] = 16'h3E01;
 buffer[323] = 16'h7B1F;
 buffer[324] = 16'h0284;
 buffer[325] = 16'h3002;
 buffer[326] = 16'h003E;
 buffer[327] = 16'h7A1C;
 buffer[328] = 16'h028A;
 buffer[329] = 16'h3E02;
 buffer[330] = 16'h003D;
 buffer[331] = 16'h7C1F;
 buffer[332] = 16'h0292;
 buffer[333] = 16'h7404;
 buffer[334] = 16'h6375;
 buffer[335] = 16'h006B;
 buffer[336] = 16'h6180;
 buffer[337] = 16'h718D;
 buffer[338] = 16'h029A;
 buffer[339] = 16'h2D04;
 buffer[340] = 16'h6F72;
 buffer[341] = 16'h0074;
 buffer[342] = 16'h6180;
 buffer[343] = 16'h6147;
 buffer[344] = 16'h6180;
 buffer[345] = 16'h6B8D;
 buffer[346] = 16'h700C;
 buffer[347] = 16'h02A6;
 buffer[348] = 16'h3202;
 buffer[349] = 16'h002F;
 buffer[350] = 16'h771C;
 buffer[351] = 16'h02B8;
 buffer[352] = 16'h3202;
 buffer[353] = 16'h002A;
 buffer[354] = 16'h751C;
 buffer[355] = 16'h02C0;
 buffer[356] = 16'h3102;
 buffer[357] = 16'h002B;
 buffer[358] = 16'h731C;
 buffer[359] = 16'h02C8;
 buffer[360] = 16'h7303;
 buffer[361] = 16'h4070;
 buffer[362] = 16'h6E81;
 buffer[363] = 16'h80FF;
 buffer[364] = 16'h730F;
 buffer[365] = 16'h02D0;
 buffer[366] = 16'h6507;
 buffer[367] = 16'h6578;
 buffer[368] = 16'h7563;
 buffer[369] = 16'h6574;
 buffer[370] = 16'h6147;
 buffer[371] = 16'h700C;
 buffer[372] = 16'h02DC;
 buffer[373] = 16'h6203;
 buffer[374] = 16'h6579;
 buffer[375] = 16'h8FFD;
 buffer[376] = 16'h6600;
 buffer[377] = 16'h6023;
 buffer[378] = 16'h710F;
 buffer[379] = 16'h02EA;
 buffer[380] = 16'h6302;
 buffer[381] = 16'h0040;
 buffer[382] = 16'h6081;
 buffer[383] = 16'h6C00;
 buffer[384] = 16'h6180;
 buffer[385] = 16'h8001;
 buffer[386] = 16'h6303;
 buffer[387] = 16'h2187;
 buffer[388] = 16'h8008;
 buffer[389] = 16'h6903;
 buffer[390] = 16'h0189;
 buffer[391] = 16'h80FF;
 buffer[392] = 16'h730F;
 buffer[393] = 16'h700C;
 buffer[394] = 16'h02F8;
 buffer[395] = 16'h6302;
 buffer[396] = 16'h0021;
 buffer[397] = 16'h6180;
 buffer[398] = 16'h80FF;
 buffer[399] = 16'h6303;
 buffer[400] = 16'h6081;
 buffer[401] = 16'h8008;
 buffer[402] = 16'h6D03;
 buffer[403] = 16'h6403;
 buffer[404] = 16'h6180;
 buffer[405] = 16'h4150;
 buffer[406] = 16'h6081;
 buffer[407] = 16'h6C00;
 buffer[408] = 16'h6180;
 buffer[409] = 16'h8001;
 buffer[410] = 16'h6303;
 buffer[411] = 16'h8000;
 buffer[412] = 16'h6703;
 buffer[413] = 16'h80FF;
 buffer[414] = 16'h6503;
 buffer[415] = 16'h6147;
 buffer[416] = 16'h6181;
 buffer[417] = 16'h6503;
 buffer[418] = 16'h6B8D;
 buffer[419] = 16'h6303;
 buffer[420] = 16'h6503;
 buffer[421] = 16'h6180;
 buffer[422] = 16'h6023;
 buffer[423] = 16'h710F;
 buffer[424] = 16'h0316;
 buffer[425] = 16'h7503;
 buffer[426] = 16'h2B6D;
 buffer[427] = 16'h6181;
 buffer[428] = 16'h6181;
 buffer[429] = 16'h6203;
 buffer[430] = 16'h6147;
 buffer[431] = 16'h6B81;
 buffer[432] = 16'h8000;
 buffer[433] = 16'h6C13;
 buffer[434] = 16'h6147;
 buffer[435] = 16'h6181;
 buffer[436] = 16'h6181;
 buffer[437] = 16'h6303;
 buffer[438] = 16'h6910;
 buffer[439] = 16'h6B8D;
 buffer[440] = 16'h6403;
 buffer[441] = 16'h6147;
 buffer[442] = 16'h6403;
 buffer[443] = 16'h6910;
 buffer[444] = 16'h6B8D;
 buffer[445] = 16'h6303;
 buffer[446] = 16'h6600;
 buffer[447] = 16'h6310;
 buffer[448] = 16'h6B8D;
 buffer[449] = 16'h718C;
 buffer[450] = 16'h0352;
 buffer[451] = 16'h6445;
 buffer[452] = 16'h766F;
 buffer[453] = 16'h7261;
 buffer[454] = 16'h6B8D;
 buffer[455] = 16'h700C;
 buffer[456] = 16'h0386;
 buffer[457] = 16'h7502;
 buffer[458] = 16'h0070;
 buffer[459] = 16'h41C6;
 buffer[460] = 16'h7E8C;
 buffer[461] = 16'h0392;
 buffer[462] = 16'h6446;
 buffer[463] = 16'h756F;
 buffer[464] = 16'h6573;
 buffer[465] = 16'h0072;
 buffer[466] = 16'h41CB;
 buffer[467] = 16'h6C00;
 buffer[468] = 16'h6B8D;
 buffer[469] = 16'h6C00;
 buffer[470] = 16'h720F;
 buffer[471] = 16'h039C;
 buffer[472] = 16'h6204;
 buffer[473] = 16'h7361;
 buffer[474] = 16'h0065;
 buffer[475] = 16'hFE80;
 buffer[476] = 16'h700C;
 buffer[477] = 16'h03B0;
 buffer[478] = 16'h7404;
 buffer[479] = 16'h6D65;
 buffer[480] = 16'h0070;
 buffer[481] = 16'hFE82;
 buffer[482] = 16'h700C;
 buffer[483] = 16'h03BC;
 buffer[484] = 16'h3E03;
 buffer[485] = 16'h6E69;
 buffer[486] = 16'hFE84;
 buffer[487] = 16'h700C;
 buffer[488] = 16'h03C8;
 buffer[489] = 16'h2304;
 buffer[490] = 16'h6974;
 buffer[491] = 16'h0062;
 buffer[492] = 16'hFE86;
 buffer[493] = 16'h700C;
 buffer[494] = 16'h03D2;
 buffer[495] = 16'h7403;
 buffer[496] = 16'h6269;
 buffer[497] = 16'hFE88;
 buffer[498] = 16'h700C;
 buffer[499] = 16'h03DE;
 buffer[500] = 16'h2705;
 buffer[501] = 16'h7665;
 buffer[502] = 16'h6C61;
 buffer[503] = 16'hFE8A;
 buffer[504] = 16'h700C;
 buffer[505] = 16'h03E8;
 buffer[506] = 16'h2706;
 buffer[507] = 16'h6261;
 buffer[508] = 16'h726F;
 buffer[509] = 16'h0074;
 buffer[510] = 16'hFE8C;
 buffer[511] = 16'h700C;
 buffer[512] = 16'h03F4;
 buffer[513] = 16'h6803;
 buffer[514] = 16'h646C;
 buffer[515] = 16'hFE8E;
 buffer[516] = 16'h700C;
 buffer[517] = 16'h0402;
 buffer[518] = 16'h6307;
 buffer[519] = 16'h6E6F;
 buffer[520] = 16'h6574;
 buffer[521] = 16'h7478;
 buffer[522] = 16'hFE90;
 buffer[523] = 16'h700C;
 buffer[524] = 16'h6413;
 buffer[525] = 16'h040C;
 buffer[526] = 16'h660E;
 buffer[527] = 16'h726F;
 buffer[528] = 16'h6874;
 buffer[529] = 16'h772D;
 buffer[530] = 16'h726F;
 buffer[531] = 16'h6C64;
 buffer[532] = 16'h7369;
 buffer[533] = 16'h0074;
 buffer[534] = 16'hFE94;
 buffer[535] = 16'h700C;
 buffer[536] = 16'h041C;
 buffer[537] = 16'h6307;
 buffer[538] = 16'h7275;
 buffer[539] = 16'h6572;
 buffer[540] = 16'h746E;
 buffer[541] = 16'hFE9A;
 buffer[542] = 16'h700C;
 buffer[543] = 16'h0432;
 buffer[544] = 16'h6402;
 buffer[545] = 16'h0070;
 buffer[546] = 16'hFE9E;
 buffer[547] = 16'h700C;
 buffer[548] = 16'h0440;
 buffer[549] = 16'h6C04;
 buffer[550] = 16'h7361;
 buffer[551] = 16'h0074;
 buffer[552] = 16'hFEA0;
 buffer[553] = 16'h700C;
 buffer[554] = 16'h044A;
 buffer[555] = 16'h2705;
 buffer[556] = 16'h6B3F;
 buffer[557] = 16'h7965;
 buffer[558] = 16'hFEA2;
 buffer[559] = 16'h700C;
 buffer[560] = 16'h0456;
 buffer[561] = 16'h2705;
 buffer[562] = 16'h6D65;
 buffer[563] = 16'h7469;
 buffer[564] = 16'hFEA4;
 buffer[565] = 16'h700C;
 buffer[566] = 16'h0462;
 buffer[567] = 16'h2705;
 buffer[568] = 16'h6F62;
 buffer[569] = 16'h746F;
 buffer[570] = 16'hFEA6;
 buffer[571] = 16'h700C;
 buffer[572] = 16'h046E;
 buffer[573] = 16'h2702;
 buffer[574] = 16'h005C;
 buffer[575] = 16'hFEA8;
 buffer[576] = 16'h700C;
 buffer[577] = 16'h047A;
 buffer[578] = 16'h2706;
 buffer[579] = 16'h616E;
 buffer[580] = 16'h656D;
 buffer[581] = 16'h003F;
 buffer[582] = 16'hFEAA;
 buffer[583] = 16'h700C;
 buffer[584] = 16'h0484;
 buffer[585] = 16'h2704;
 buffer[586] = 16'h2C24;
 buffer[587] = 16'h006E;
 buffer[588] = 16'hFEAC;
 buffer[589] = 16'h700C;
 buffer[590] = 16'h0492;
 buffer[591] = 16'h2706;
 buffer[592] = 16'h766F;
 buffer[593] = 16'h7265;
 buffer[594] = 16'h0074;
 buffer[595] = 16'hFEAE;
 buffer[596] = 16'h700C;
 buffer[597] = 16'h049E;
 buffer[598] = 16'h2702;
 buffer[599] = 16'h003B;
 buffer[600] = 16'hFEB0;
 buffer[601] = 16'h700C;
 buffer[602] = 16'h04AC;
 buffer[603] = 16'h2707;
 buffer[604] = 16'h7263;
 buffer[605] = 16'h6165;
 buffer[606] = 16'h6574;
 buffer[607] = 16'hFEB2;
 buffer[608] = 16'h700C;
 buffer[609] = 16'h04B6;
 buffer[610] = 16'h6402;
 buffer[611] = 16'h0021;
 buffer[612] = 16'h6180;
 buffer[613] = 16'h6181;
 buffer[614] = 16'h6023;
 buffer[615] = 16'h6103;
 buffer[616] = 16'h6310;
 buffer[617] = 16'h6023;
 buffer[618] = 16'h710F;
 buffer[619] = 16'h04C4;
 buffer[620] = 16'h6402;
 buffer[621] = 16'h0040;
 buffer[622] = 16'h6081;
 buffer[623] = 16'h6310;
 buffer[624] = 16'h6C00;
 buffer[625] = 16'h6180;
 buffer[626] = 16'h7C0C;
 buffer[627] = 16'h04D8;
 buffer[628] = 16'h3F04;
 buffer[629] = 16'h7564;
 buffer[630] = 16'h0070;
 buffer[631] = 16'h6081;
 buffer[632] = 16'h227A;
 buffer[633] = 16'h708D;
 buffer[634] = 16'h700C;
 buffer[635] = 16'h04E8;
 buffer[636] = 16'h7203;
 buffer[637] = 16'h746F;
 buffer[638] = 16'h6147;
 buffer[639] = 16'h6180;
 buffer[640] = 16'h6B8D;
 buffer[641] = 16'h718C;
 buffer[642] = 16'h04F8;
 buffer[643] = 16'h3205;
 buffer[644] = 16'h7264;
 buffer[645] = 16'h706F;
 buffer[646] = 16'h6103;
 buffer[647] = 16'h710F;
 buffer[648] = 16'h0506;
 buffer[649] = 16'h3204;
 buffer[650] = 16'h7564;
 buffer[651] = 16'h0070;
 buffer[652] = 16'h6181;
 buffer[653] = 16'h718D;
 buffer[654] = 16'h0512;
 buffer[655] = 16'h6E06;
 buffer[656] = 16'h6765;
 buffer[657] = 16'h7461;
 buffer[658] = 16'h0065;
 buffer[659] = 16'h761C;
 buffer[660] = 16'h051E;
 buffer[661] = 16'h6407;
 buffer[662] = 16'h656E;
 buffer[663] = 16'h6167;
 buffer[664] = 16'h6574;
 buffer[665] = 16'h805F;
 buffer[666] = 16'h6600;
 buffer[667] = 16'h4264;
 buffer[668] = 16'h8053;
 buffer[669] = 16'h6600;
 buffer[670] = 16'h026E;
 buffer[671] = 16'h052A;
 buffer[672] = 16'h2D01;
 buffer[673] = 16'h781F;
 buffer[674] = 16'h0540;
 buffer[675] = 16'h6103;
 buffer[676] = 16'h7362;
 buffer[677] = 16'h7D1C;
 buffer[678] = 16'h0546;
 buffer[679] = 16'h6D03;
 buffer[680] = 16'h7861;
 buffer[681] = 16'h7E1F;
 buffer[682] = 16'h054E;
 buffer[683] = 16'h6D03;
 buffer[684] = 16'h6E69;
 buffer[685] = 16'h7F1F;
 buffer[686] = 16'h0556;
 buffer[687] = 16'h7706;
 buffer[688] = 16'h7469;
 buffer[689] = 16'h6968;
 buffer[690] = 16'h006E;
 buffer[691] = 16'h6181;
 buffer[692] = 16'h42A1;
 buffer[693] = 16'h6147;
 buffer[694] = 16'h42A1;
 buffer[695] = 16'h6B8D;
 buffer[696] = 16'h7F0F;
 buffer[697] = 16'h055E;
 buffer[698] = 16'h6D03;
 buffer[699] = 16'h212F;
 buffer[700] = 16'h802D;
 buffer[701] = 16'h6600;
 buffer[702] = 16'h6023;
 buffer[703] = 16'h6103;
 buffer[704] = 16'h802F;
 buffer[705] = 16'h6600;
 buffer[706] = 16'h0264;
 buffer[707] = 16'h0574;
 buffer[708] = 16'h6D03;
 buffer[709] = 16'h3F2F;
 buffer[710] = 16'h802C;
 buffer[711] = 16'h6600;
 buffer[712] = 16'h6023;
 buffer[713] = 16'h6103;
 buffer[714] = 16'h802C;
 buffer[715] = 16'h6600;
 buffer[716] = 16'h6C00;
 buffer[717] = 16'h6010;
 buffer[718] = 16'h22CA;
 buffer[719] = 16'h802E;
 buffer[720] = 16'h6600;
 buffer[721] = 16'h6C00;
 buffer[722] = 16'h802F;
 buffer[723] = 16'h6600;
 buffer[724] = 16'h7C0C;
 buffer[725] = 16'h0588;
 buffer[726] = 16'h7506;
 buffer[727] = 16'h2F6D;
 buffer[728] = 16'h6F6D;
 buffer[729] = 16'h0064;
 buffer[730] = 16'h42BC;
 buffer[731] = 16'h8001;
 buffer[732] = 16'h02C6;
 buffer[733] = 16'h05AC;
 buffer[734] = 16'h6D05;
 buffer[735] = 16'h6D2F;
 buffer[736] = 16'h646F;
 buffer[737] = 16'h42BC;
 buffer[738] = 16'h8002;
 buffer[739] = 16'h02C6;
 buffer[740] = 16'h05BC;
 buffer[741] = 16'h2F02;
 buffer[742] = 16'h0021;
 buffer[743] = 16'h802A;
 buffer[744] = 16'h6600;
 buffer[745] = 16'h6023;
 buffer[746] = 16'h6103;
 buffer[747] = 16'h802B;
 buffer[748] = 16'h6600;
 buffer[749] = 16'h6023;
 buffer[750] = 16'h6103;
 buffer[751] = 16'h8001;
 buffer[752] = 16'h8029;
 buffer[753] = 16'h6600;
 buffer[754] = 16'h6023;
 buffer[755] = 16'h710F;
 buffer[756] = 16'h05CA;
 buffer[757] = 16'h2F04;
 buffer[758] = 16'h6F6D;
 buffer[759] = 16'h0064;
 buffer[760] = 16'h42E7;
 buffer[761] = 16'h8029;
 buffer[762] = 16'h6600;
 buffer[763] = 16'h6C00;
 buffer[764] = 16'h6010;
 buffer[765] = 16'h22F9;
 buffer[766] = 16'h802A;
 buffer[767] = 16'h6600;
 buffer[768] = 16'h6C00;
 buffer[769] = 16'h802B;
 buffer[770] = 16'h6600;
 buffer[771] = 16'h7C0C;
 buffer[772] = 16'h05EA;
 buffer[773] = 16'h6D03;
 buffer[774] = 16'h646F;
 buffer[775] = 16'h42F8;
 buffer[776] = 16'h710F;
 buffer[777] = 16'h060A;
 buffer[778] = 16'h2F01;
 buffer[779] = 16'h42F8;
 buffer[780] = 16'h700F;
 buffer[781] = 16'h0614;
 buffer[782] = 16'h6D03;
 buffer[783] = 16'h212A;
 buffer[784] = 16'h8028;
 buffer[785] = 16'h6600;
 buffer[786] = 16'h6023;
 buffer[787] = 16'h6103;
 buffer[788] = 16'h8027;
 buffer[789] = 16'h6600;
 buffer[790] = 16'h6023;
 buffer[791] = 16'h710F;
 buffer[792] = 16'h061C;
 buffer[793] = 16'h6D03;
 buffer[794] = 16'h3F2A;
 buffer[795] = 16'h8026;
 buffer[796] = 16'h6600;
 buffer[797] = 16'h6023;
 buffer[798] = 16'h6103;
 buffer[799] = 16'h8028;
 buffer[800] = 16'h6600;
 buffer[801] = 16'h026E;
 buffer[802] = 16'h0632;
 buffer[803] = 16'h7503;
 buffer[804] = 16'h2A6D;
 buffer[805] = 16'h4310;
 buffer[806] = 16'h8001;
 buffer[807] = 16'h031B;
 buffer[808] = 16'h0646;
 buffer[809] = 16'h6D02;
 buffer[810] = 16'h002A;
 buffer[811] = 16'h4310;
 buffer[812] = 16'h8002;
 buffer[813] = 16'h031B;
 buffer[814] = 16'h0652;
 buffer[815] = 16'h2A01;
 buffer[816] = 16'h741F;
 buffer[817] = 16'h065E;
 buffer[818] = 16'h2A05;
 buffer[819] = 16'h6D2F;
 buffer[820] = 16'h646F;
 buffer[821] = 16'h6147;
 buffer[822] = 16'h432B;
 buffer[823] = 16'h6B8D;
 buffer[824] = 16'h02E1;
 buffer[825] = 16'h0664;
 buffer[826] = 16'h2A02;
 buffer[827] = 16'h002F;
 buffer[828] = 16'h4335;
 buffer[829] = 16'h700F;
 buffer[830] = 16'h0674;
 buffer[831] = 16'h6305;
 buffer[832] = 16'h6C65;
 buffer[833] = 16'h2B6C;
 buffer[834] = 16'h8002;
 buffer[835] = 16'h720F;
 buffer[836] = 16'h067E;
 buffer[837] = 16'h6305;
 buffer[838] = 16'h6C65;
 buffer[839] = 16'h2D6C;
 buffer[840] = 16'h8002;
 buffer[841] = 16'h02A1;
 buffer[842] = 16'h068A;
 buffer[843] = 16'h6305;
 buffer[844] = 16'h6C65;
 buffer[845] = 16'h736C;
 buffer[846] = 16'h8001;
 buffer[847] = 16'h7D0F;
 buffer[848] = 16'h0696;
 buffer[849] = 16'h6202;
 buffer[850] = 16'h006C;
 buffer[851] = 16'h8020;
 buffer[852] = 16'h700C;
 buffer[853] = 16'h06A2;
 buffer[854] = 16'h3E05;
 buffer[855] = 16'h6863;
 buffer[856] = 16'h7261;
 buffer[857] = 16'h807F;
 buffer[858] = 16'h6303;
 buffer[859] = 16'h6081;
 buffer[860] = 16'h807F;
 buffer[861] = 16'h4353;
 buffer[862] = 16'h42B3;
 buffer[863] = 16'h2362;
 buffer[864] = 16'h6103;
 buffer[865] = 16'h805F;
 buffer[866] = 16'h700C;
 buffer[867] = 16'h700C;
 buffer[868] = 16'h06AC;
 buffer[869] = 16'h2B02;
 buffer[870] = 16'h0021;
 buffer[871] = 16'h4150;
 buffer[872] = 16'h6C00;
 buffer[873] = 16'h6203;
 buffer[874] = 16'h6180;
 buffer[875] = 16'h6023;
 buffer[876] = 16'h710F;
 buffer[877] = 16'h06CA;
 buffer[878] = 16'h3202;
 buffer[879] = 16'h0021;
 buffer[880] = 16'h6180;
 buffer[881] = 16'h6181;
 buffer[882] = 16'h6023;
 buffer[883] = 16'h6103;
 buffer[884] = 16'h4342;
 buffer[885] = 16'h6023;
 buffer[886] = 16'h710F;
 buffer[887] = 16'h06DC;
 buffer[888] = 16'h3202;
 buffer[889] = 16'h0040;
 buffer[890] = 16'h6081;
 buffer[891] = 16'h4342;
 buffer[892] = 16'h6C00;
 buffer[893] = 16'h6180;
 buffer[894] = 16'h7C0C;
 buffer[895] = 16'h06F0;
 buffer[896] = 16'h6305;
 buffer[897] = 16'h756F;
 buffer[898] = 16'h746E;
 buffer[899] = 16'h6081;
 buffer[900] = 16'h6310;
 buffer[901] = 16'h6180;
 buffer[902] = 16'h017E;
 buffer[903] = 16'h0700;
 buffer[904] = 16'h6804;
 buffer[905] = 16'h7265;
 buffer[906] = 16'h0065;
 buffer[907] = 16'hFE9E;
 buffer[908] = 16'h7C0C;
 buffer[909] = 16'h0710;
 buffer[910] = 16'h6107;
 buffer[911] = 16'h696C;
 buffer[912] = 16'h6E67;
 buffer[913] = 16'h6465;
 buffer[914] = 16'h6081;
 buffer[915] = 16'h8000;
 buffer[916] = 16'h8002;
 buffer[917] = 16'h42DA;
 buffer[918] = 16'h6103;
 buffer[919] = 16'h6081;
 buffer[920] = 16'h239C;
 buffer[921] = 16'h8002;
 buffer[922] = 16'h6180;
 buffer[923] = 16'h42A1;
 buffer[924] = 16'h720F;
 buffer[925] = 16'h071C;
 buffer[926] = 16'h6105;
 buffer[927] = 16'h696C;
 buffer[928] = 16'h6E67;
 buffer[929] = 16'h438B;
 buffer[930] = 16'h4392;
 buffer[931] = 16'hFE9E;
 buffer[932] = 16'h6023;
 buffer[933] = 16'h710F;
 buffer[934] = 16'h073C;
 buffer[935] = 16'h7003;
 buffer[936] = 16'h6461;
 buffer[937] = 16'h438B;
 buffer[938] = 16'h8050;
 buffer[939] = 16'h6203;
 buffer[940] = 16'h0392;
 buffer[941] = 16'h074E;
 buffer[942] = 16'h4008;
 buffer[943] = 16'h7865;
 buffer[944] = 16'h6365;
 buffer[945] = 16'h7475;
 buffer[946] = 16'h0065;
 buffer[947] = 16'h6C00;
 buffer[948] = 16'h4277;
 buffer[949] = 16'h23B7;
 buffer[950] = 16'h0172;
 buffer[951] = 16'h700C;
 buffer[952] = 16'h075C;
 buffer[953] = 16'h6604;
 buffer[954] = 16'h6C69;
 buffer[955] = 16'h006C;
 buffer[956] = 16'h6180;
 buffer[957] = 16'h6147;
 buffer[958] = 16'h6180;
 buffer[959] = 16'h03C3;
 buffer[960] = 16'h428C;
 buffer[961] = 16'h418D;
 buffer[962] = 16'h6310;
 buffer[963] = 16'h6B81;
 buffer[964] = 16'h23C9;
 buffer[965] = 16'h6B8D;
 buffer[966] = 16'h6A00;
 buffer[967] = 16'h6147;
 buffer[968] = 16'h03C0;
 buffer[969] = 16'h6B8D;
 buffer[970] = 16'h6103;
 buffer[971] = 16'h0286;
 buffer[972] = 16'h0772;
 buffer[973] = 16'h6505;
 buffer[974] = 16'h6172;
 buffer[975] = 16'h6573;
 buffer[976] = 16'h8000;
 buffer[977] = 16'h03BC;
 buffer[978] = 16'h079A;
 buffer[979] = 16'h6405;
 buffer[980] = 16'h6769;
 buffer[981] = 16'h7469;
 buffer[982] = 16'h8009;
 buffer[983] = 16'h6181;
 buffer[984] = 16'h6803;
 buffer[985] = 16'h8007;
 buffer[986] = 16'h6303;
 buffer[987] = 16'h6203;
 buffer[988] = 16'h8030;
 buffer[989] = 16'h720F;
 buffer[990] = 16'h07A6;
 buffer[991] = 16'h6507;
 buffer[992] = 16'h7478;
 buffer[993] = 16'h6172;
 buffer[994] = 16'h7463;
 buffer[995] = 16'h8000;
 buffer[996] = 16'h6180;
 buffer[997] = 16'h42DA;
 buffer[998] = 16'h6180;
 buffer[999] = 16'h03D6;
 buffer[1000] = 16'h07BE;
 buffer[1001] = 16'h3C02;
 buffer[1002] = 16'h0023;
 buffer[1003] = 16'h43A9;
 buffer[1004] = 16'hFE8E;
 buffer[1005] = 16'h6023;
 buffer[1006] = 16'h710F;
 buffer[1007] = 16'h07D2;
 buffer[1008] = 16'h6804;
 buffer[1009] = 16'h6C6F;
 buffer[1010] = 16'h0064;
 buffer[1011] = 16'hFE8E;
 buffer[1012] = 16'h6C00;
 buffer[1013] = 16'h6A00;
 buffer[1014] = 16'h6081;
 buffer[1015] = 16'hFE8E;
 buffer[1016] = 16'h6023;
 buffer[1017] = 16'h6103;
 buffer[1018] = 16'h018D;
 buffer[1019] = 16'h07E0;
 buffer[1020] = 16'h2301;
 buffer[1021] = 16'hFE80;
 buffer[1022] = 16'h6C00;
 buffer[1023] = 16'h43E3;
 buffer[1024] = 16'h03F3;
 buffer[1025] = 16'h07F8;
 buffer[1026] = 16'h2302;
 buffer[1027] = 16'h0073;
 buffer[1028] = 16'h43FD;
 buffer[1029] = 16'h6081;
 buffer[1030] = 16'h2408;
 buffer[1031] = 16'h0404;
 buffer[1032] = 16'h700C;
 buffer[1033] = 16'h0804;
 buffer[1034] = 16'h7304;
 buffer[1035] = 16'h6769;
 buffer[1036] = 16'h006E;
 buffer[1037] = 16'h6910;
 buffer[1038] = 16'h2411;
 buffer[1039] = 16'h802D;
 buffer[1040] = 16'h03F3;
 buffer[1041] = 16'h700C;
 buffer[1042] = 16'h0814;
 buffer[1043] = 16'h2302;
 buffer[1044] = 16'h003E;
 buffer[1045] = 16'h6103;
 buffer[1046] = 16'hFE8E;
 buffer[1047] = 16'h6C00;
 buffer[1048] = 16'h43A9;
 buffer[1049] = 16'h6181;
 buffer[1050] = 16'h02A1;
 buffer[1051] = 16'h0826;
 buffer[1052] = 16'h7303;
 buffer[1053] = 16'h7274;
 buffer[1054] = 16'h6081;
 buffer[1055] = 16'h6147;
 buffer[1056] = 16'h6D10;
 buffer[1057] = 16'h43EB;
 buffer[1058] = 16'h4404;
 buffer[1059] = 16'h6B8D;
 buffer[1060] = 16'h440D;
 buffer[1061] = 16'h0415;
 buffer[1062] = 16'h0838;
 buffer[1063] = 16'h6803;
 buffer[1064] = 16'h7865;
 buffer[1065] = 16'h8010;
 buffer[1066] = 16'hFE80;
 buffer[1067] = 16'h6023;
 buffer[1068] = 16'h710F;
 buffer[1069] = 16'h084E;
 buffer[1070] = 16'h6407;
 buffer[1071] = 16'h6365;
 buffer[1072] = 16'h6D69;
 buffer[1073] = 16'h6C61;
 buffer[1074] = 16'h800A;
 buffer[1075] = 16'hFE80;
 buffer[1076] = 16'h6023;
 buffer[1077] = 16'h710F;
 buffer[1078] = 16'h085C;
 buffer[1079] = 16'h6406;
 buffer[1080] = 16'h6769;
 buffer[1081] = 16'h7469;
 buffer[1082] = 16'h003F;
 buffer[1083] = 16'h6147;
 buffer[1084] = 16'h8030;
 buffer[1085] = 16'h42A1;
 buffer[1086] = 16'h8009;
 buffer[1087] = 16'h6181;
 buffer[1088] = 16'h6803;
 buffer[1089] = 16'h244E;
 buffer[1090] = 16'h6081;
 buffer[1091] = 16'h8020;
 buffer[1092] = 16'h6B13;
 buffer[1093] = 16'h2448;
 buffer[1094] = 16'h8020;
 buffer[1095] = 16'h42A1;
 buffer[1096] = 16'h8007;
 buffer[1097] = 16'h42A1;
 buffer[1098] = 16'h6081;
 buffer[1099] = 16'h800A;
 buffer[1100] = 16'h6803;
 buffer[1101] = 16'h6403;
 buffer[1102] = 16'h6081;
 buffer[1103] = 16'h6B8D;
 buffer[1104] = 16'h7F0F;
 buffer[1105] = 16'h086E;
 buffer[1106] = 16'h6E07;
 buffer[1107] = 16'h6D75;
 buffer[1108] = 16'h6562;
 buffer[1109] = 16'h3F72;
 buffer[1110] = 16'hFE80;
 buffer[1111] = 16'h6C00;
 buffer[1112] = 16'h6147;
 buffer[1113] = 16'h8000;
 buffer[1114] = 16'h6181;
 buffer[1115] = 16'h4383;
 buffer[1116] = 16'h6181;
 buffer[1117] = 16'h417E;
 buffer[1118] = 16'h8024;
 buffer[1119] = 16'h6703;
 buffer[1120] = 16'h2466;
 buffer[1121] = 16'h4429;
 buffer[1122] = 16'h6180;
 buffer[1123] = 16'h6310;
 buffer[1124] = 16'h6180;
 buffer[1125] = 16'h6A00;
 buffer[1126] = 16'h6181;
 buffer[1127] = 16'h417E;
 buffer[1128] = 16'h802D;
 buffer[1129] = 16'h6703;
 buffer[1130] = 16'h6147;
 buffer[1131] = 16'h6180;
 buffer[1132] = 16'h6B81;
 buffer[1133] = 16'h42A1;
 buffer[1134] = 16'h6180;
 buffer[1135] = 16'h6B81;
 buffer[1136] = 16'h6203;
 buffer[1137] = 16'h4277;
 buffer[1138] = 16'h2497;
 buffer[1139] = 16'h6A00;
 buffer[1140] = 16'h6147;
 buffer[1141] = 16'h6081;
 buffer[1142] = 16'h6147;
 buffer[1143] = 16'h417E;
 buffer[1144] = 16'hFE80;
 buffer[1145] = 16'h6C00;
 buffer[1146] = 16'h443B;
 buffer[1147] = 16'h2491;
 buffer[1148] = 16'h6180;
 buffer[1149] = 16'hFE80;
 buffer[1150] = 16'h6C00;
 buffer[1151] = 16'h6413;
 buffer[1152] = 16'h6203;
 buffer[1153] = 16'h6B8D;
 buffer[1154] = 16'h6310;
 buffer[1155] = 16'h6B81;
 buffer[1156] = 16'h2489;
 buffer[1157] = 16'h6B8D;
 buffer[1158] = 16'h6A00;
 buffer[1159] = 16'h6147;
 buffer[1160] = 16'h0475;
 buffer[1161] = 16'h6B8D;
 buffer[1162] = 16'h6103;
 buffer[1163] = 16'h6B81;
 buffer[1164] = 16'h6003;
 buffer[1165] = 16'h248F;
 buffer[1166] = 16'h6610;
 buffer[1167] = 16'h6180;
 buffer[1168] = 16'h0496;
 buffer[1169] = 16'h6B8D;
 buffer[1170] = 16'h6B8D;
 buffer[1171] = 16'h4286;
 buffer[1172] = 16'h4286;
 buffer[1173] = 16'h8000;
 buffer[1174] = 16'h6081;
 buffer[1175] = 16'h6B8D;
 buffer[1176] = 16'h4286;
 buffer[1177] = 16'h6B8D;
 buffer[1178] = 16'hFE80;
 buffer[1179] = 16'h6023;
 buffer[1180] = 16'h710F;
 buffer[1181] = 16'h08A4;
 buffer[1182] = 16'h3F03;
 buffer[1183] = 16'h7872;
 buffer[1184] = 16'h8FFE;
 buffer[1185] = 16'h6600;
 buffer[1186] = 16'h6C00;
 buffer[1187] = 16'h8001;
 buffer[1188] = 16'h6303;
 buffer[1189] = 16'h711C;
 buffer[1190] = 16'h093C;
 buffer[1191] = 16'h7403;
 buffer[1192] = 16'h2178;
 buffer[1193] = 16'h8FFE;
 buffer[1194] = 16'h6600;
 buffer[1195] = 16'h6C00;
 buffer[1196] = 16'h8002;
 buffer[1197] = 16'h6303;
 buffer[1198] = 16'h6010;
 buffer[1199] = 16'h24A9;
 buffer[1200] = 16'h6081;
 buffer[1201] = 16'h8FFF;
 buffer[1202] = 16'h6600;
 buffer[1203] = 16'h6023;
 buffer[1204] = 16'h6103;
 buffer[1205] = 16'h80DF;
 buffer[1206] = 16'h6600;
 buffer[1207] = 16'h6C00;
 buffer[1208] = 16'h6010;
 buffer[1209] = 16'h24B5;
 buffer[1210] = 16'h80DF;
 buffer[1211] = 16'h6600;
 buffer[1212] = 16'h6023;
 buffer[1213] = 16'h710F;
 buffer[1214] = 16'h094E;
 buffer[1215] = 16'h3F04;
 buffer[1216] = 16'h656B;
 buffer[1217] = 16'h0079;
 buffer[1218] = 16'hFEA2;
 buffer[1219] = 16'h03B3;
 buffer[1220] = 16'h097E;
 buffer[1221] = 16'h6504;
 buffer[1222] = 16'h696D;
 buffer[1223] = 16'h0074;
 buffer[1224] = 16'hFEA4;
 buffer[1225] = 16'h03B3;
 buffer[1226] = 16'h098A;
 buffer[1227] = 16'h6B03;
 buffer[1228] = 16'h7965;
 buffer[1229] = 16'h44C2;
 buffer[1230] = 16'h24CD;
 buffer[1231] = 16'h8FFF;
 buffer[1232] = 16'h6600;
 buffer[1233] = 16'h7C0C;
 buffer[1234] = 16'h0996;
 buffer[1235] = 16'h6E04;
 buffer[1236] = 16'h6675;
 buffer[1237] = 16'h003F;
 buffer[1238] = 16'h44C2;
 buffer[1239] = 16'h6081;
 buffer[1240] = 16'h24DD;
 buffer[1241] = 16'h6103;
 buffer[1242] = 16'h44CD;
 buffer[1243] = 16'h800D;
 buffer[1244] = 16'h770F;
 buffer[1245] = 16'h700C;
 buffer[1246] = 16'h09A6;
 buffer[1247] = 16'h7305;
 buffer[1248] = 16'h6170;
 buffer[1249] = 16'h6563;
 buffer[1250] = 16'h4353;
 buffer[1251] = 16'h04C8;
 buffer[1252] = 16'h09BE;
 buffer[1253] = 16'h7306;
 buffer[1254] = 16'h6170;
 buffer[1255] = 16'h6563;
 buffer[1256] = 16'h0073;
 buffer[1257] = 16'h8000;
 buffer[1258] = 16'h6E13;
 buffer[1259] = 16'h6147;
 buffer[1260] = 16'h04EE;
 buffer[1261] = 16'h44E2;
 buffer[1262] = 16'h6B81;
 buffer[1263] = 16'h24F4;
 buffer[1264] = 16'h6B8D;
 buffer[1265] = 16'h6A00;
 buffer[1266] = 16'h6147;
 buffer[1267] = 16'h04ED;
 buffer[1268] = 16'h6B8D;
 buffer[1269] = 16'h710F;
 buffer[1270] = 16'h09CA;
 buffer[1271] = 16'h7404;
 buffer[1272] = 16'h7079;
 buffer[1273] = 16'h0065;
 buffer[1274] = 16'h6147;
 buffer[1275] = 16'h04FE;
 buffer[1276] = 16'h4383;
 buffer[1277] = 16'h44C8;
 buffer[1278] = 16'h6B81;
 buffer[1279] = 16'h2504;
 buffer[1280] = 16'h6B8D;
 buffer[1281] = 16'h6A00;
 buffer[1282] = 16'h6147;
 buffer[1283] = 16'h04FC;
 buffer[1284] = 16'h6B8D;
 buffer[1285] = 16'h6103;
 buffer[1286] = 16'h710F;
 buffer[1287] = 16'h09EE;
 buffer[1288] = 16'h6302;
 buffer[1289] = 16'h0072;
 buffer[1290] = 16'h800D;
 buffer[1291] = 16'h44C8;
 buffer[1292] = 16'h800A;
 buffer[1293] = 16'h04C8;
 buffer[1294] = 16'h0A10;
 buffer[1295] = 16'h6443;
 buffer[1296] = 16'h246F;
 buffer[1297] = 16'h6B8D;
 buffer[1298] = 16'h6B81;
 buffer[1299] = 16'h6B8D;
 buffer[1300] = 16'h4383;
 buffer[1301] = 16'h6203;
 buffer[1302] = 16'h4392;
 buffer[1303] = 16'h6147;
 buffer[1304] = 16'h6180;
 buffer[1305] = 16'h6147;
 buffer[1306] = 16'h700C;
 buffer[1307] = 16'h0A1E;
 buffer[1308] = 16'h2443;
 buffer[1309] = 16'h7C22;
 buffer[1310] = 16'h4511;
 buffer[1311] = 16'h700C;
 buffer[1312] = 16'h0A38;
 buffer[1313] = 16'h2E02;
 buffer[1314] = 16'h0024;
 buffer[1315] = 16'h4383;
 buffer[1316] = 16'h04FA;
 buffer[1317] = 16'h0A42;
 buffer[1318] = 16'h2E43;
 buffer[1319] = 16'h7C22;
 buffer[1320] = 16'h4511;
 buffer[1321] = 16'h0523;
 buffer[1322] = 16'h0A4C;
 buffer[1323] = 16'h2E02;
 buffer[1324] = 16'h0072;
 buffer[1325] = 16'h6147;
 buffer[1326] = 16'h441E;
 buffer[1327] = 16'h6B8D;
 buffer[1328] = 16'h6181;
 buffer[1329] = 16'h42A1;
 buffer[1330] = 16'h44E9;
 buffer[1331] = 16'h04FA;
 buffer[1332] = 16'h0A56;
 buffer[1333] = 16'h7503;
 buffer[1334] = 16'h722E;
 buffer[1335] = 16'h6147;
 buffer[1336] = 16'h43EB;
 buffer[1337] = 16'h4404;
 buffer[1338] = 16'h4415;
 buffer[1339] = 16'h6B8D;
 buffer[1340] = 16'h6181;
 buffer[1341] = 16'h42A1;
 buffer[1342] = 16'h44E9;
 buffer[1343] = 16'h04FA;
 buffer[1344] = 16'h0A6A;
 buffer[1345] = 16'h7502;
 buffer[1346] = 16'h002E;
 buffer[1347] = 16'h43EB;
 buffer[1348] = 16'h4404;
 buffer[1349] = 16'h4415;
 buffer[1350] = 16'h44E2;
 buffer[1351] = 16'h04FA;
 buffer[1352] = 16'h0A82;
 buffer[1353] = 16'h2E01;
 buffer[1354] = 16'hFE80;
 buffer[1355] = 16'h6C00;
 buffer[1356] = 16'h800A;
 buffer[1357] = 16'h6503;
 buffer[1358] = 16'h2550;
 buffer[1359] = 16'h0543;
 buffer[1360] = 16'h441E;
 buffer[1361] = 16'h44E2;
 buffer[1362] = 16'h04FA;
 buffer[1363] = 16'h0A92;
 buffer[1364] = 16'h6305;
 buffer[1365] = 16'h6F6D;
 buffer[1366] = 16'h6576;
 buffer[1367] = 16'h6147;
 buffer[1368] = 16'h0561;
 buffer[1369] = 16'h6147;
 buffer[1370] = 16'h6081;
 buffer[1371] = 16'h417E;
 buffer[1372] = 16'h6B81;
 buffer[1373] = 16'h418D;
 buffer[1374] = 16'h6310;
 buffer[1375] = 16'h6B8D;
 buffer[1376] = 16'h6310;
 buffer[1377] = 16'h6B81;
 buffer[1378] = 16'h2567;
 buffer[1379] = 16'h6B8D;
 buffer[1380] = 16'h6A00;
 buffer[1381] = 16'h6147;
 buffer[1382] = 16'h0559;
 buffer[1383] = 16'h6B8D;
 buffer[1384] = 16'h6103;
 buffer[1385] = 16'h0286;
 buffer[1386] = 16'h0AA8;
 buffer[1387] = 16'h7005;
 buffer[1388] = 16'h6361;
 buffer[1389] = 16'h246B;
 buffer[1390] = 16'h6081;
 buffer[1391] = 16'h6147;
 buffer[1392] = 16'h428C;
 buffer[1393] = 16'h6023;
 buffer[1394] = 16'h6103;
 buffer[1395] = 16'h6310;
 buffer[1396] = 16'h6180;
 buffer[1397] = 16'h4557;
 buffer[1398] = 16'h6B8D;
 buffer[1399] = 16'h700C;
 buffer[1400] = 16'h0AD6;
 buffer[1401] = 16'h3F01;
 buffer[1402] = 16'h6C00;
 buffer[1403] = 16'h054A;
 buffer[1404] = 16'h0AF2;
 buffer[1405] = 16'h2807;
 buffer[1406] = 16'h6170;
 buffer[1407] = 16'h7372;
 buffer[1408] = 16'h2965;
 buffer[1409] = 16'hFE82;
 buffer[1410] = 16'h6023;
 buffer[1411] = 16'h6103;
 buffer[1412] = 16'h6181;
 buffer[1413] = 16'h6147;
 buffer[1414] = 16'h6081;
 buffer[1415] = 16'h25CC;
 buffer[1416] = 16'h6A00;
 buffer[1417] = 16'hFE82;
 buffer[1418] = 16'h6C00;
 buffer[1419] = 16'h4353;
 buffer[1420] = 16'h6703;
 buffer[1421] = 16'h25A8;
 buffer[1422] = 16'h6147;
 buffer[1423] = 16'h4383;
 buffer[1424] = 16'hFE82;
 buffer[1425] = 16'h6C00;
 buffer[1426] = 16'h6180;
 buffer[1427] = 16'h42A1;
 buffer[1428] = 16'h6910;
 buffer[1429] = 16'h6600;
 buffer[1430] = 16'h6B81;
 buffer[1431] = 16'h6A10;
 buffer[1432] = 16'h6303;
 buffer[1433] = 16'h25A6;
 buffer[1434] = 16'h6B81;
 buffer[1435] = 16'h25A0;
 buffer[1436] = 16'h6B8D;
 buffer[1437] = 16'h6A00;
 buffer[1438] = 16'h6147;
 buffer[1439] = 16'h058F;
 buffer[1440] = 16'h6B8D;
 buffer[1441] = 16'h6103;
 buffer[1442] = 16'h6B8D;
 buffer[1443] = 16'h6103;
 buffer[1444] = 16'h8000;
 buffer[1445] = 16'h708D;
 buffer[1446] = 16'h6A00;
 buffer[1447] = 16'h6B8D;
 buffer[1448] = 16'h6181;
 buffer[1449] = 16'h6180;
 buffer[1450] = 16'h6147;
 buffer[1451] = 16'h4383;
 buffer[1452] = 16'hFE82;
 buffer[1453] = 16'h6C00;
 buffer[1454] = 16'h6180;
 buffer[1455] = 16'h42A1;
 buffer[1456] = 16'hFE82;
 buffer[1457] = 16'h6C00;
 buffer[1458] = 16'h4353;
 buffer[1459] = 16'h6703;
 buffer[1460] = 16'h25B6;
 buffer[1461] = 16'h6910;
 buffer[1462] = 16'h25C2;
 buffer[1463] = 16'h6B81;
 buffer[1464] = 16'h25BD;
 buffer[1465] = 16'h6B8D;
 buffer[1466] = 16'h6A00;
 buffer[1467] = 16'h6147;
 buffer[1468] = 16'h05AB;
 buffer[1469] = 16'h6B8D;
 buffer[1470] = 16'h6103;
 buffer[1471] = 16'h6081;
 buffer[1472] = 16'h6147;
 buffer[1473] = 16'h05C7;
 buffer[1474] = 16'h6B8D;
 buffer[1475] = 16'h6103;
 buffer[1476] = 16'h6081;
 buffer[1477] = 16'h6147;
 buffer[1478] = 16'h6A00;
 buffer[1479] = 16'h6181;
 buffer[1480] = 16'h42A1;
 buffer[1481] = 16'h6B8D;
 buffer[1482] = 16'h6B8D;
 buffer[1483] = 16'h02A1;
 buffer[1484] = 16'h6181;
 buffer[1485] = 16'h6B8D;
 buffer[1486] = 16'h02A1;
 buffer[1487] = 16'h0AFA;
 buffer[1488] = 16'h7005;
 buffer[1489] = 16'h7261;
 buffer[1490] = 16'h6573;
 buffer[1491] = 16'h6147;
 buffer[1492] = 16'hFE88;
 buffer[1493] = 16'h6C00;
 buffer[1494] = 16'hFE84;
 buffer[1495] = 16'h6C00;
 buffer[1496] = 16'h6203;
 buffer[1497] = 16'hFE86;
 buffer[1498] = 16'h6C00;
 buffer[1499] = 16'hFE84;
 buffer[1500] = 16'h6C00;
 buffer[1501] = 16'h42A1;
 buffer[1502] = 16'h6B8D;
 buffer[1503] = 16'h4581;
 buffer[1504] = 16'hFE84;
 buffer[1505] = 16'h0367;
 buffer[1506] = 16'h0BA0;
 buffer[1507] = 16'h2E82;
 buffer[1508] = 16'h0028;
 buffer[1509] = 16'h8029;
 buffer[1510] = 16'h45D3;
 buffer[1511] = 16'h04FA;
 buffer[1512] = 16'h0BC6;
 buffer[1513] = 16'h2881;
 buffer[1514] = 16'h8029;
 buffer[1515] = 16'h45D3;
 buffer[1516] = 16'h0286;
 buffer[1517] = 16'h0BD2;
 buffer[1518] = 16'h3C83;
 buffer[1519] = 16'h3E5C;
 buffer[1520] = 16'hFE86;
 buffer[1521] = 16'h6C00;
 buffer[1522] = 16'hFE84;
 buffer[1523] = 16'h6023;
 buffer[1524] = 16'h710F;
 buffer[1525] = 16'h0BDC;
 buffer[1526] = 16'h5C81;
 buffer[1527] = 16'hFEA8;
 buffer[1528] = 16'h03B3;
 buffer[1529] = 16'h0BEC;
 buffer[1530] = 16'h7704;
 buffer[1531] = 16'h726F;
 buffer[1532] = 16'h0064;
 buffer[1533] = 16'h45D3;
 buffer[1534] = 16'h438B;
 buffer[1535] = 16'h4342;
 buffer[1536] = 16'h056E;
 buffer[1537] = 16'h0BF4;
 buffer[1538] = 16'h7405;
 buffer[1539] = 16'h6B6F;
 buffer[1540] = 16'h6E65;
 buffer[1541] = 16'h4353;
 buffer[1542] = 16'h05FD;
 buffer[1543] = 16'h0C04;
 buffer[1544] = 16'h6E05;
 buffer[1545] = 16'h6D61;
 buffer[1546] = 16'h3E65;
 buffer[1547] = 16'h4383;
 buffer[1548] = 16'h801F;
 buffer[1549] = 16'h6303;
 buffer[1550] = 16'h6203;
 buffer[1551] = 16'h0392;
 buffer[1552] = 16'h0C10;
 buffer[1553] = 16'h7305;
 buffer[1554] = 16'h6D61;
 buffer[1555] = 16'h3F65;
 buffer[1556] = 16'h6A00;
 buffer[1557] = 16'h6147;
 buffer[1558] = 16'h0624;
 buffer[1559] = 16'h6181;
 buffer[1560] = 16'h6B81;
 buffer[1561] = 16'h6203;
 buffer[1562] = 16'h417E;
 buffer[1563] = 16'h6181;
 buffer[1564] = 16'h6B81;
 buffer[1565] = 16'h6203;
 buffer[1566] = 16'h417E;
 buffer[1567] = 16'h42A1;
 buffer[1568] = 16'h4277;
 buffer[1569] = 16'h2624;
 buffer[1570] = 16'h6B8D;
 buffer[1571] = 16'h710F;
 buffer[1572] = 16'h6B81;
 buffer[1573] = 16'h262A;
 buffer[1574] = 16'h6B8D;
 buffer[1575] = 16'h6A00;
 buffer[1576] = 16'h6147;
 buffer[1577] = 16'h0617;
 buffer[1578] = 16'h6B8D;
 buffer[1579] = 16'h6103;
 buffer[1580] = 16'h8000;
 buffer[1581] = 16'h700C;
 buffer[1582] = 16'h0C22;
 buffer[1583] = 16'h6604;
 buffer[1584] = 16'h6E69;
 buffer[1585] = 16'h0064;
 buffer[1586] = 16'h6180;
 buffer[1587] = 16'h6081;
 buffer[1588] = 16'h417E;
 buffer[1589] = 16'hFE82;
 buffer[1590] = 16'h6023;
 buffer[1591] = 16'h6103;
 buffer[1592] = 16'h6081;
 buffer[1593] = 16'h6C00;
 buffer[1594] = 16'h6147;
 buffer[1595] = 16'h4342;
 buffer[1596] = 16'h6180;
 buffer[1597] = 16'h6C00;
 buffer[1598] = 16'h6081;
 buffer[1599] = 16'h2650;
 buffer[1600] = 16'h6081;
 buffer[1601] = 16'h6C00;
 buffer[1602] = 16'hFF1F;
 buffer[1603] = 16'h6303;
 buffer[1604] = 16'h6B81;
 buffer[1605] = 16'h6503;
 buffer[1606] = 16'h264B;
 buffer[1607] = 16'h4342;
 buffer[1608] = 16'h8000;
 buffer[1609] = 16'h6600;
 buffer[1610] = 16'h064F;
 buffer[1611] = 16'h4342;
 buffer[1612] = 16'hFE82;
 buffer[1613] = 16'h6C00;
 buffer[1614] = 16'h4614;
 buffer[1615] = 16'h0655;
 buffer[1616] = 16'h6B8D;
 buffer[1617] = 16'h6103;
 buffer[1618] = 16'h6180;
 buffer[1619] = 16'h4348;
 buffer[1620] = 16'h718C;
 buffer[1621] = 16'h265A;
 buffer[1622] = 16'h8002;
 buffer[1623] = 16'h434E;
 buffer[1624] = 16'h42A1;
 buffer[1625] = 16'h063D;
 buffer[1626] = 16'h6B8D;
 buffer[1627] = 16'h6103;
 buffer[1628] = 16'h6003;
 buffer[1629] = 16'h4348;
 buffer[1630] = 16'h6081;
 buffer[1631] = 16'h460B;
 buffer[1632] = 16'h718C;
 buffer[1633] = 16'h0C5E;
 buffer[1634] = 16'h3C07;
 buffer[1635] = 16'h616E;
 buffer[1636] = 16'h656D;
 buffer[1637] = 16'h3E3F;
 buffer[1638] = 16'hFE90;
 buffer[1639] = 16'h6081;
 buffer[1640] = 16'h437A;
 buffer[1641] = 16'h6503;
 buffer[1642] = 16'h266C;
 buffer[1643] = 16'h4348;
 buffer[1644] = 16'h6147;
 buffer[1645] = 16'h6B8D;
 buffer[1646] = 16'h4342;
 buffer[1647] = 16'h6081;
 buffer[1648] = 16'h6147;
 buffer[1649] = 16'h6C00;
 buffer[1650] = 16'h4277;
 buffer[1651] = 16'h2679;
 buffer[1652] = 16'h4632;
 buffer[1653] = 16'h4277;
 buffer[1654] = 16'h266D;
 buffer[1655] = 16'h6B8D;
 buffer[1656] = 16'h710F;
 buffer[1657] = 16'h6B8D;
 buffer[1658] = 16'h6103;
 buffer[1659] = 16'h8000;
 buffer[1660] = 16'h700C;
 buffer[1661] = 16'h0CC4;
 buffer[1662] = 16'h6E05;
 buffer[1663] = 16'h6D61;
 buffer[1664] = 16'h3F65;
 buffer[1665] = 16'hFEAA;
 buffer[1666] = 16'h03B3;
 buffer[1667] = 16'h0CFC;
 buffer[1668] = 16'h5E02;
 buffer[1669] = 16'h0068;
 buffer[1670] = 16'h6147;
 buffer[1671] = 16'h6181;
 buffer[1672] = 16'h6B81;
 buffer[1673] = 16'h6803;
 buffer[1674] = 16'h6081;
 buffer[1675] = 16'h2691;
 buffer[1676] = 16'h8008;
 buffer[1677] = 16'h6081;
 buffer[1678] = 16'h44C8;
 buffer[1679] = 16'h44E2;
 buffer[1680] = 16'h44C8;
 buffer[1681] = 16'h6B8D;
 buffer[1682] = 16'h720F;
 buffer[1683] = 16'h0D08;
 buffer[1684] = 16'h7403;
 buffer[1685] = 16'h7061;
 buffer[1686] = 16'h6081;
 buffer[1687] = 16'h44C8;
 buffer[1688] = 16'h6181;
 buffer[1689] = 16'h418D;
 buffer[1690] = 16'h731C;
 buffer[1691] = 16'h0D28;
 buffer[1692] = 16'h6B04;
 buffer[1693] = 16'h6174;
 buffer[1694] = 16'h0070;
 buffer[1695] = 16'h6081;
 buffer[1696] = 16'h800D;
 buffer[1697] = 16'h6503;
 buffer[1698] = 16'h26A9;
 buffer[1699] = 16'h8008;
 buffer[1700] = 16'h6503;
 buffer[1701] = 16'h26A8;
 buffer[1702] = 16'h4353;
 buffer[1703] = 16'h0696;
 buffer[1704] = 16'h0686;
 buffer[1705] = 16'h6103;
 buffer[1706] = 16'h6003;
 buffer[1707] = 16'h708D;
 buffer[1708] = 16'h0D38;
 buffer[1709] = 16'h6106;
 buffer[1710] = 16'h6363;
 buffer[1711] = 16'h7065;
 buffer[1712] = 16'h0074;
 buffer[1713] = 16'h6181;
 buffer[1714] = 16'h6203;
 buffer[1715] = 16'h6181;
 buffer[1716] = 16'h428C;
 buffer[1717] = 16'h6503;
 buffer[1718] = 16'h26C2;
 buffer[1719] = 16'h44CD;
 buffer[1720] = 16'h6081;
 buffer[1721] = 16'h4353;
 buffer[1722] = 16'h42A1;
 buffer[1723] = 16'h807F;
 buffer[1724] = 16'h6F03;
 buffer[1725] = 16'h26C0;
 buffer[1726] = 16'h4696;
 buffer[1727] = 16'h06C1;
 buffer[1728] = 16'h469F;
 buffer[1729] = 16'h06B4;
 buffer[1730] = 16'h6103;
 buffer[1731] = 16'h6181;
 buffer[1732] = 16'h02A1;
 buffer[1733] = 16'h0D5A;
 buffer[1734] = 16'h7105;
 buffer[1735] = 16'h6575;
 buffer[1736] = 16'h7972;
 buffer[1737] = 16'hFE88;
 buffer[1738] = 16'h6C00;
 buffer[1739] = 16'h8050;
 buffer[1740] = 16'h46B1;
 buffer[1741] = 16'hFE86;
 buffer[1742] = 16'h6023;
 buffer[1743] = 16'h6103;
 buffer[1744] = 16'h6103;
 buffer[1745] = 16'h8000;
 buffer[1746] = 16'hFE84;
 buffer[1747] = 16'h6023;
 buffer[1748] = 16'h710F;
 buffer[1749] = 16'h0D8C;
 buffer[1750] = 16'h6106;
 buffer[1751] = 16'h6F62;
 buffer[1752] = 16'h7472;
 buffer[1753] = 16'h0032;
 buffer[1754] = 16'h4511;
 buffer[1755] = 16'h710F;
 buffer[1756] = 16'h0DAC;
 buffer[1757] = 16'h6106;
 buffer[1758] = 16'h6F62;
 buffer[1759] = 16'h7472;
 buffer[1760] = 16'h0031;
 buffer[1761] = 16'h44E2;
 buffer[1762] = 16'h4523;
 buffer[1763] = 16'h803F;
 buffer[1764] = 16'h44C8;
 buffer[1765] = 16'h450A;
 buffer[1766] = 16'hFE8C;
 buffer[1767] = 16'h43B3;
 buffer[1768] = 16'h06DA;
 buffer[1769] = 16'h0DBA;
 buffer[1770] = 16'h3C49;
 buffer[1771] = 16'h613F;
 buffer[1772] = 16'h6F62;
 buffer[1773] = 16'h7472;
 buffer[1774] = 16'h3E22;
 buffer[1775] = 16'h26F2;
 buffer[1776] = 16'h4511;
 buffer[1777] = 16'h06E1;
 buffer[1778] = 16'h06DA;
 buffer[1779] = 16'h0DD4;
 buffer[1780] = 16'h6606;
 buffer[1781] = 16'h726F;
 buffer[1782] = 16'h6567;
 buffer[1783] = 16'h0074;
 buffer[1784] = 16'h4605;
 buffer[1785] = 16'h4681;
 buffer[1786] = 16'h4277;
 buffer[1787] = 16'h270A;
 buffer[1788] = 16'h4348;
 buffer[1789] = 16'h6081;
 buffer[1790] = 16'hFE9E;
 buffer[1791] = 16'h6023;
 buffer[1792] = 16'h6103;
 buffer[1793] = 16'h6C00;
 buffer[1794] = 16'h6081;
 buffer[1795] = 16'hFE90;
 buffer[1796] = 16'h6023;
 buffer[1797] = 16'h6103;
 buffer[1798] = 16'hFEA0;
 buffer[1799] = 16'h6023;
 buffer[1800] = 16'h6103;
 buffer[1801] = 16'h710F;
 buffer[1802] = 16'h06E1;
 buffer[1803] = 16'h0DE8;
 buffer[1804] = 16'h240A;
 buffer[1805] = 16'h6E69;
 buffer[1806] = 16'h6574;
 buffer[1807] = 16'h7072;
 buffer[1808] = 16'h6572;
 buffer[1809] = 16'h0074;
 buffer[1810] = 16'h4681;
 buffer[1811] = 16'h4277;
 buffer[1812] = 16'h2722;
 buffer[1813] = 16'h6C00;
 buffer[1814] = 16'h8040;
 buffer[1815] = 16'h6303;
 buffer[1816] = 16'h46EF;
 buffer[1817] = 16'h630C;
 buffer[1818] = 16'h6D6F;
 buffer[1819] = 16'h6970;
 buffer[1820] = 16'h656C;
 buffer[1821] = 16'h6F2D;
 buffer[1822] = 16'h6C6E;
 buffer[1823] = 16'h0079;
 buffer[1824] = 16'h0172;
 buffer[1825] = 16'h0726;
 buffer[1826] = 16'h4456;
 buffer[1827] = 16'h2725;
 buffer[1828] = 16'h700C;
 buffer[1829] = 16'h06E1;
 buffer[1830] = 16'h0E18;
 buffer[1831] = 16'h5B81;
 buffer[1832] = 16'h8E24;
 buffer[1833] = 16'hFE8A;
 buffer[1834] = 16'h6023;
 buffer[1835] = 16'h710F;
 buffer[1836] = 16'h0E4E;
 buffer[1837] = 16'h2E03;
 buffer[1838] = 16'h6B6F;
 buffer[1839] = 16'h8E24;
 buffer[1840] = 16'hFE8A;
 buffer[1841] = 16'h6C00;
 buffer[1842] = 16'h6703;
 buffer[1843] = 16'h2737;
 buffer[1844] = 16'h4528;
 buffer[1845] = 16'h2003;
 buffer[1846] = 16'h6B6F;
 buffer[1847] = 16'h050A;
 buffer[1848] = 16'h0E5A;
 buffer[1849] = 16'h6504;
 buffer[1850] = 16'h6176;
 buffer[1851] = 16'h006C;
 buffer[1852] = 16'h4605;
 buffer[1853] = 16'h6081;
 buffer[1854] = 16'h417E;
 buffer[1855] = 16'h2743;
 buffer[1856] = 16'hFE8A;
 buffer[1857] = 16'h43B3;
 buffer[1858] = 16'h073C;
 buffer[1859] = 16'h6103;
 buffer[1860] = 16'h072F;
 buffer[1861] = 16'h0E72;
 buffer[1862] = 16'h2445;
 buffer[1863] = 16'h7665;
 buffer[1864] = 16'h6C61;
 buffer[1865] = 16'hFE84;
 buffer[1866] = 16'h6C00;
 buffer[1867] = 16'h6147;
 buffer[1868] = 16'hFE86;
 buffer[1869] = 16'h6C00;
 buffer[1870] = 16'h6147;
 buffer[1871] = 16'hFE88;
 buffer[1872] = 16'h6C00;
 buffer[1873] = 16'h6147;
 buffer[1874] = 16'hFE84;
 buffer[1875] = 16'h8000;
 buffer[1876] = 16'h6180;
 buffer[1877] = 16'h6023;
 buffer[1878] = 16'h6103;
 buffer[1879] = 16'hFE86;
 buffer[1880] = 16'h6023;
 buffer[1881] = 16'h6103;
 buffer[1882] = 16'hFE88;
 buffer[1883] = 16'h6023;
 buffer[1884] = 16'h6103;
 buffer[1885] = 16'h473C;
 buffer[1886] = 16'h6B8D;
 buffer[1887] = 16'hFE88;
 buffer[1888] = 16'h6023;
 buffer[1889] = 16'h6103;
 buffer[1890] = 16'h6B8D;
 buffer[1891] = 16'hFE86;
 buffer[1892] = 16'h6023;
 buffer[1893] = 16'h6103;
 buffer[1894] = 16'h6B8D;
 buffer[1895] = 16'hFE84;
 buffer[1896] = 16'h6023;
 buffer[1897] = 16'h710F;
 buffer[1898] = 16'h0E8C;
 buffer[1899] = 16'h7006;
 buffer[1900] = 16'h6572;
 buffer[1901] = 16'h6573;
 buffer[1902] = 16'h0074;
 buffer[1903] = 16'hFF00;
 buffer[1904] = 16'hFE86;
 buffer[1905] = 16'h4342;
 buffer[1906] = 16'h6023;
 buffer[1907] = 16'h710F;
 buffer[1908] = 16'h0ED6;
 buffer[1909] = 16'h7104;
 buffer[1910] = 16'h6975;
 buffer[1911] = 16'h0074;
 buffer[1912] = 16'h4728;
 buffer[1913] = 16'h46C9;
 buffer[1914] = 16'h473C;
 buffer[1915] = 16'h0779;
 buffer[1916] = 16'h700C;
 buffer[1917] = 16'h0EEA;
 buffer[1918] = 16'h6105;
 buffer[1919] = 16'h6F62;
 buffer[1920] = 16'h7472;
 buffer[1921] = 16'h6103;
 buffer[1922] = 16'h476F;
 buffer[1923] = 16'h472F;
 buffer[1924] = 16'h0778;
 buffer[1925] = 16'h0EFC;
 buffer[1926] = 16'h2701;
 buffer[1927] = 16'h4605;
 buffer[1928] = 16'h4681;
 buffer[1929] = 16'h278B;
 buffer[1930] = 16'h700C;
 buffer[1931] = 16'h06E1;
 buffer[1932] = 16'h0F0C;
 buffer[1933] = 16'h6105;
 buffer[1934] = 16'h6C6C;
 buffer[1935] = 16'h746F;
 buffer[1936] = 16'h4392;
 buffer[1937] = 16'hFE9E;
 buffer[1938] = 16'h0367;
 buffer[1939] = 16'h0F1A;
 buffer[1940] = 16'h2C01;
 buffer[1941] = 16'h438B;
 buffer[1942] = 16'h6081;
 buffer[1943] = 16'h4342;
 buffer[1944] = 16'hFE9E;
 buffer[1945] = 16'h6023;
 buffer[1946] = 16'h6103;
 buffer[1947] = 16'h6023;
 buffer[1948] = 16'h710F;
 buffer[1949] = 16'h0F28;
 buffer[1950] = 16'h6345;
 buffer[1951] = 16'h6C61;
 buffer[1952] = 16'h2C6C;
 buffer[1953] = 16'h8001;
 buffer[1954] = 16'h6903;
 buffer[1955] = 16'hC000;
 buffer[1956] = 16'h6403;
 buffer[1957] = 16'h0795;
 buffer[1958] = 16'h0F3C;
 buffer[1959] = 16'h3F47;
 buffer[1960] = 16'h7262;
 buffer[1961] = 16'h6E61;
 buffer[1962] = 16'h6863;
 buffer[1963] = 16'h8001;
 buffer[1964] = 16'h6903;
 buffer[1965] = 16'hA000;
 buffer[1966] = 16'h6403;
 buffer[1967] = 16'h0795;
 buffer[1968] = 16'h0F4E;
 buffer[1969] = 16'h6246;
 buffer[1970] = 16'h6172;
 buffer[1971] = 16'h636E;
 buffer[1972] = 16'h0068;
 buffer[1973] = 16'h8001;
 buffer[1974] = 16'h6903;
 buffer[1975] = 16'h8000;
 buffer[1976] = 16'h6403;
 buffer[1977] = 16'h0795;
 buffer[1978] = 16'h0F62;
 buffer[1979] = 16'h5B89;
 buffer[1980] = 16'h6F63;
 buffer[1981] = 16'h706D;
 buffer[1982] = 16'h6C69;
 buffer[1983] = 16'h5D65;
 buffer[1984] = 16'h4787;
 buffer[1985] = 16'h07A1;
 buffer[1986] = 16'h0F76;
 buffer[1987] = 16'h6347;
 buffer[1988] = 16'h6D6F;
 buffer[1989] = 16'h6970;
 buffer[1990] = 16'h656C;
 buffer[1991] = 16'h6B8D;
 buffer[1992] = 16'h6081;
 buffer[1993] = 16'h6C00;
 buffer[1994] = 16'h4795;
 buffer[1995] = 16'h4342;
 buffer[1996] = 16'h6147;
 buffer[1997] = 16'h700C;
 buffer[1998] = 16'h0F86;
 buffer[1999] = 16'h7287;
 buffer[2000] = 16'h6365;
 buffer[2001] = 16'h7275;
 buffer[2002] = 16'h6573;
 buffer[2003] = 16'hFEA0;
 buffer[2004] = 16'h6C00;
 buffer[2005] = 16'h460B;
 buffer[2006] = 16'h07A1;
 buffer[2007] = 16'h0F9E;
 buffer[2008] = 16'h7004;
 buffer[2009] = 16'h6369;
 buffer[2010] = 16'h006B;
 buffer[2011] = 16'h6081;
 buffer[2012] = 16'h6510;
 buffer[2013] = 16'h6510;
 buffer[2014] = 16'h80C0;
 buffer[2015] = 16'h6203;
 buffer[2016] = 16'h6147;
 buffer[2017] = 16'h700C;
 buffer[2018] = 16'h0FB0;
 buffer[2019] = 16'h6C87;
 buffer[2020] = 16'h7469;
 buffer[2021] = 16'h7265;
 buffer[2022] = 16'h6C61;
 buffer[2023] = 16'h6081;
 buffer[2024] = 16'hFFFF;
 buffer[2025] = 16'h6600;
 buffer[2026] = 16'h6303;
 buffer[2027] = 16'h27F3;
 buffer[2028] = 16'h8000;
 buffer[2029] = 16'h6600;
 buffer[2030] = 16'h6503;
 buffer[2031] = 16'h47E7;
 buffer[2032] = 16'h47C7;
 buffer[2033] = 16'h6600;
 buffer[2034] = 16'h07F7;
 buffer[2035] = 16'hFFFF;
 buffer[2036] = 16'h6600;
 buffer[2037] = 16'h6403;
 buffer[2038] = 16'h0795;
 buffer[2039] = 16'h700C;
 buffer[2040] = 16'h0FC6;
 buffer[2041] = 16'h5B83;
 buffer[2042] = 16'h5D27;
 buffer[2043] = 16'h4787;
 buffer[2044] = 16'h07E7;
 buffer[2045] = 16'h0FF2;
 buffer[2046] = 16'h2403;
 buffer[2047] = 16'h222C;
 buffer[2048] = 16'h8022;
 buffer[2049] = 16'h45D3;
 buffer[2050] = 16'h438B;
 buffer[2051] = 16'h456E;
 buffer[2052] = 16'h4383;
 buffer[2053] = 16'h6203;
 buffer[2054] = 16'h4392;
 buffer[2055] = 16'hFE9E;
 buffer[2056] = 16'h6023;
 buffer[2057] = 16'h710F;
 buffer[2058] = 16'h0FFC;
 buffer[2059] = 16'h66C3;
 buffer[2060] = 16'h726F;
 buffer[2061] = 16'h47C7;
 buffer[2062] = 16'h4113;
 buffer[2063] = 16'h038B;
 buffer[2064] = 16'h1016;
 buffer[2065] = 16'h62C5;
 buffer[2066] = 16'h6765;
 buffer[2067] = 16'h6E69;
 buffer[2068] = 16'h038B;
 buffer[2069] = 16'h1022;
 buffer[2070] = 16'h2846;
 buffer[2071] = 16'h656E;
 buffer[2072] = 16'h7478;
 buffer[2073] = 16'h0029;
 buffer[2074] = 16'h6B8D;
 buffer[2075] = 16'h6B8D;
 buffer[2076] = 16'h4277;
 buffer[2077] = 16'h2823;
 buffer[2078] = 16'h6A00;
 buffer[2079] = 16'h6147;
 buffer[2080] = 16'h6C00;
 buffer[2081] = 16'h6147;
 buffer[2082] = 16'h700C;
 buffer[2083] = 16'h4342;
 buffer[2084] = 16'h6147;
 buffer[2085] = 16'h700C;
 buffer[2086] = 16'h102C;
 buffer[2087] = 16'h6EC4;
 buffer[2088] = 16'h7865;
 buffer[2089] = 16'h0074;
 buffer[2090] = 16'h47C7;
 buffer[2091] = 16'h481A;
 buffer[2092] = 16'h0795;
 buffer[2093] = 16'h104E;
 buffer[2094] = 16'h2844;
 buffer[2095] = 16'h6F64;
 buffer[2096] = 16'h0029;
 buffer[2097] = 16'h6B8D;
 buffer[2098] = 16'h6081;
 buffer[2099] = 16'h6147;
 buffer[2100] = 16'h6180;
 buffer[2101] = 16'h427E;
 buffer[2102] = 16'h6147;
 buffer[2103] = 16'h6147;
 buffer[2104] = 16'h4342;
 buffer[2105] = 16'h6147;
 buffer[2106] = 16'h700C;
 buffer[2107] = 16'h105C;
 buffer[2108] = 16'h64C2;
 buffer[2109] = 16'h006F;
 buffer[2110] = 16'h47C7;
 buffer[2111] = 16'h4831;
 buffer[2112] = 16'h8000;
 buffer[2113] = 16'h4795;
 buffer[2114] = 16'h038B;
 buffer[2115] = 16'h1078;
 buffer[2116] = 16'h2847;
 buffer[2117] = 16'h656C;
 buffer[2118] = 16'h7661;
 buffer[2119] = 16'h2965;
 buffer[2120] = 16'h6B8D;
 buffer[2121] = 16'h6103;
 buffer[2122] = 16'h6B8D;
 buffer[2123] = 16'h6103;
 buffer[2124] = 16'h6B8D;
 buffer[2125] = 16'h710F;
 buffer[2126] = 16'h1088;
 buffer[2127] = 16'h6CC5;
 buffer[2128] = 16'h6165;
 buffer[2129] = 16'h6576;
 buffer[2130] = 16'h47C7;
 buffer[2131] = 16'h4848;
 buffer[2132] = 16'h700C;
 buffer[2133] = 16'h109E;
 buffer[2134] = 16'h2846;
 buffer[2135] = 16'h6F6C;
 buffer[2136] = 16'h706F;
 buffer[2137] = 16'h0029;
 buffer[2138] = 16'h6B8D;
 buffer[2139] = 16'h6B8D;
 buffer[2140] = 16'h6310;
 buffer[2141] = 16'h6B8D;
 buffer[2142] = 16'h428C;
 buffer[2143] = 16'h6213;
 buffer[2144] = 16'h2866;
 buffer[2145] = 16'h6147;
 buffer[2146] = 16'h6147;
 buffer[2147] = 16'h6C00;
 buffer[2148] = 16'h6147;
 buffer[2149] = 16'h700C;
 buffer[2150] = 16'h6147;
 buffer[2151] = 16'h6A00;
 buffer[2152] = 16'h6147;
 buffer[2153] = 16'h4342;
 buffer[2154] = 16'h6147;
 buffer[2155] = 16'h700C;
 buffer[2156] = 16'h10AC;
 buffer[2157] = 16'h2848;
 buffer[2158] = 16'h6E75;
 buffer[2159] = 16'h6F6C;
 buffer[2160] = 16'h706F;
 buffer[2161] = 16'h0029;
 buffer[2162] = 16'h6B8D;
 buffer[2163] = 16'h6B8D;
 buffer[2164] = 16'h6103;
 buffer[2165] = 16'h6B8D;
 buffer[2166] = 16'h6103;
 buffer[2167] = 16'h6B8D;
 buffer[2168] = 16'h6103;
 buffer[2169] = 16'h6147;
 buffer[2170] = 16'h700C;
 buffer[2171] = 16'h10DA;
 buffer[2172] = 16'h75C6;
 buffer[2173] = 16'h6C6E;
 buffer[2174] = 16'h6F6F;
 buffer[2175] = 16'h0070;
 buffer[2176] = 16'h47C7;
 buffer[2177] = 16'h4872;
 buffer[2178] = 16'h700C;
 buffer[2179] = 16'h10F8;
 buffer[2180] = 16'h2845;
 buffer[2181] = 16'h643F;
 buffer[2182] = 16'h296F;
 buffer[2183] = 16'h428C;
 buffer[2184] = 16'h6213;
 buffer[2185] = 16'h2894;
 buffer[2186] = 16'h6B8D;
 buffer[2187] = 16'h6081;
 buffer[2188] = 16'h6147;
 buffer[2189] = 16'h6180;
 buffer[2190] = 16'h427E;
 buffer[2191] = 16'h6147;
 buffer[2192] = 16'h6147;
 buffer[2193] = 16'h4342;
 buffer[2194] = 16'h6147;
 buffer[2195] = 16'h700C;
 buffer[2196] = 16'h0286;
 buffer[2197] = 16'h700C;
 buffer[2198] = 16'h1108;
 buffer[2199] = 16'h3FC3;
 buffer[2200] = 16'h6F64;
 buffer[2201] = 16'h47C7;
 buffer[2202] = 16'h4887;
 buffer[2203] = 16'h8000;
 buffer[2204] = 16'h4795;
 buffer[2205] = 16'h038B;
 buffer[2206] = 16'h112E;
 buffer[2207] = 16'h6CC4;
 buffer[2208] = 16'h6F6F;
 buffer[2209] = 16'h0070;
 buffer[2210] = 16'h47C7;
 buffer[2211] = 16'h485A;
 buffer[2212] = 16'h6081;
 buffer[2213] = 16'h4795;
 buffer[2214] = 16'h47C7;
 buffer[2215] = 16'h4872;
 buffer[2216] = 16'h4348;
 buffer[2217] = 16'h438B;
 buffer[2218] = 16'h8001;
 buffer[2219] = 16'h6903;
 buffer[2220] = 16'h6180;
 buffer[2221] = 16'h6023;
 buffer[2222] = 16'h710F;
 buffer[2223] = 16'h113E;
 buffer[2224] = 16'h2847;
 buffer[2225] = 16'h6C2B;
 buffer[2226] = 16'h6F6F;
 buffer[2227] = 16'h2970;
 buffer[2228] = 16'h6B8D;
 buffer[2229] = 16'h6180;
 buffer[2230] = 16'h6B8D;
 buffer[2231] = 16'h6B8D;
 buffer[2232] = 16'h428C;
 buffer[2233] = 16'h42A1;
 buffer[2234] = 16'h6147;
 buffer[2235] = 16'h8002;
 buffer[2236] = 16'h47DB;
 buffer[2237] = 16'h6B81;
 buffer[2238] = 16'h6203;
 buffer[2239] = 16'h6B81;
 buffer[2240] = 16'h6503;
 buffer[2241] = 16'h6910;
 buffer[2242] = 16'h6010;
 buffer[2243] = 16'h8003;
 buffer[2244] = 16'h47DB;
 buffer[2245] = 16'h6B8D;
 buffer[2246] = 16'h6503;
 buffer[2247] = 16'h6910;
 buffer[2248] = 16'h6010;
 buffer[2249] = 16'h6403;
 buffer[2250] = 16'h28D1;
 buffer[2251] = 16'h6147;
 buffer[2252] = 16'h6203;
 buffer[2253] = 16'h6147;
 buffer[2254] = 16'h6C00;
 buffer[2255] = 16'h6147;
 buffer[2256] = 16'h700C;
 buffer[2257] = 16'h6147;
 buffer[2258] = 16'h6147;
 buffer[2259] = 16'h6103;
 buffer[2260] = 16'h4342;
 buffer[2261] = 16'h6147;
 buffer[2262] = 16'h700C;
 buffer[2263] = 16'h1160;
 buffer[2264] = 16'h2BC5;
 buffer[2265] = 16'h6F6C;
 buffer[2266] = 16'h706F;
 buffer[2267] = 16'h47C7;
 buffer[2268] = 16'h48B4;
 buffer[2269] = 16'h6081;
 buffer[2270] = 16'h4795;
 buffer[2271] = 16'h47C7;
 buffer[2272] = 16'h4872;
 buffer[2273] = 16'h4348;
 buffer[2274] = 16'h438B;
 buffer[2275] = 16'h8001;
 buffer[2276] = 16'h6903;
 buffer[2277] = 16'h6180;
 buffer[2278] = 16'h6023;
 buffer[2279] = 16'h710F;
 buffer[2280] = 16'h11B0;
 buffer[2281] = 16'h2843;
 buffer[2282] = 16'h2969;
 buffer[2283] = 16'h6B8D;
 buffer[2284] = 16'h6B8D;
 buffer[2285] = 16'h4150;
 buffer[2286] = 16'h6147;
 buffer[2287] = 16'h6147;
 buffer[2288] = 16'h700C;
 buffer[2289] = 16'h11D2;
 buffer[2290] = 16'h69C1;
 buffer[2291] = 16'h47C7;
 buffer[2292] = 16'h48EB;
 buffer[2293] = 16'h700C;
 buffer[2294] = 16'h11E4;
 buffer[2295] = 16'h75C5;
 buffer[2296] = 16'h746E;
 buffer[2297] = 16'h6C69;
 buffer[2298] = 16'h07AB;
 buffer[2299] = 16'h11EE;
 buffer[2300] = 16'h61C5;
 buffer[2301] = 16'h6167;
 buffer[2302] = 16'h6E69;
 buffer[2303] = 16'h07B5;
 buffer[2304] = 16'h11F8;
 buffer[2305] = 16'h69C2;
 buffer[2306] = 16'h0066;
 buffer[2307] = 16'h438B;
 buffer[2308] = 16'h8000;
 buffer[2309] = 16'h07AB;
 buffer[2310] = 16'h1202;
 buffer[2311] = 16'h74C4;
 buffer[2312] = 16'h6568;
 buffer[2313] = 16'h006E;
 buffer[2314] = 16'h438B;
 buffer[2315] = 16'h8001;
 buffer[2316] = 16'h6903;
 buffer[2317] = 16'h6181;
 buffer[2318] = 16'h6C00;
 buffer[2319] = 16'h6403;
 buffer[2320] = 16'h6180;
 buffer[2321] = 16'h6023;
 buffer[2322] = 16'h710F;
 buffer[2323] = 16'h120E;
 buffer[2324] = 16'h72C6;
 buffer[2325] = 16'h7065;
 buffer[2326] = 16'h6165;
 buffer[2327] = 16'h0074;
 buffer[2328] = 16'h47B5;
 buffer[2329] = 16'h090A;
 buffer[2330] = 16'h1228;
 buffer[2331] = 16'h73C4;
 buffer[2332] = 16'h696B;
 buffer[2333] = 16'h0070;
 buffer[2334] = 16'h438B;
 buffer[2335] = 16'h8000;
 buffer[2336] = 16'h07B5;
 buffer[2337] = 16'h1236;
 buffer[2338] = 16'h61C3;
 buffer[2339] = 16'h7466;
 buffer[2340] = 16'h6103;
 buffer[2341] = 16'h491E;
 buffer[2342] = 16'h4814;
 buffer[2343] = 16'h718C;
 buffer[2344] = 16'h1244;
 buffer[2345] = 16'h65C4;
 buffer[2346] = 16'h736C;
 buffer[2347] = 16'h0065;
 buffer[2348] = 16'h491E;
 buffer[2349] = 16'h6180;
 buffer[2350] = 16'h090A;
 buffer[2351] = 16'h1252;
 buffer[2352] = 16'h77C5;
 buffer[2353] = 16'h6968;
 buffer[2354] = 16'h656C;
 buffer[2355] = 16'h4903;
 buffer[2356] = 16'h718C;
 buffer[2357] = 16'h1260;
 buffer[2358] = 16'h2846;
 buffer[2359] = 16'h6163;
 buffer[2360] = 16'h6573;
 buffer[2361] = 16'h0029;
 buffer[2362] = 16'h6B8D;
 buffer[2363] = 16'h6180;
 buffer[2364] = 16'h6147;
 buffer[2365] = 16'h6147;
 buffer[2366] = 16'h700C;
 buffer[2367] = 16'h126C;
 buffer[2368] = 16'h63C4;
 buffer[2369] = 16'h7361;
 buffer[2370] = 16'h0065;
 buffer[2371] = 16'h47C7;
 buffer[2372] = 16'h493A;
 buffer[2373] = 16'h8030;
 buffer[2374] = 16'h700C;
 buffer[2375] = 16'h1280;
 buffer[2376] = 16'h2844;
 buffer[2377] = 16'h666F;
 buffer[2378] = 16'h0029;
 buffer[2379] = 16'h6B8D;
 buffer[2380] = 16'h6B81;
 buffer[2381] = 16'h6180;
 buffer[2382] = 16'h6147;
 buffer[2383] = 16'h770F;
 buffer[2384] = 16'h1290;
 buffer[2385] = 16'h6FC2;
 buffer[2386] = 16'h0066;
 buffer[2387] = 16'h47C7;
 buffer[2388] = 16'h494B;
 buffer[2389] = 16'h0903;
 buffer[2390] = 16'h12A2;
 buffer[2391] = 16'h65C5;
 buffer[2392] = 16'h646E;
 buffer[2393] = 16'h666F;
 buffer[2394] = 16'h492C;
 buffer[2395] = 16'h8031;
 buffer[2396] = 16'h700C;
 buffer[2397] = 16'h12AE;
 buffer[2398] = 16'h2809;
 buffer[2399] = 16'h6E65;
 buffer[2400] = 16'h6364;
 buffer[2401] = 16'h7361;
 buffer[2402] = 16'h2965;
 buffer[2403] = 16'h6B8D;
 buffer[2404] = 16'h6B8D;
 buffer[2405] = 16'h6103;
 buffer[2406] = 16'h6147;
 buffer[2407] = 16'h700C;
 buffer[2408] = 16'h12BC;
 buffer[2409] = 16'h65C7;
 buffer[2410] = 16'h646E;
 buffer[2411] = 16'h6163;
 buffer[2412] = 16'h6573;
 buffer[2413] = 16'h6081;
 buffer[2414] = 16'h8031;
 buffer[2415] = 16'h6703;
 buffer[2416] = 16'h2974;
 buffer[2417] = 16'h6103;
 buffer[2418] = 16'h490A;
 buffer[2419] = 16'h096D;
 buffer[2420] = 16'h8030;
 buffer[2421] = 16'h6213;
 buffer[2422] = 16'h46EF;
 buffer[2423] = 16'h6213;
 buffer[2424] = 16'h6461;
 buffer[2425] = 16'h6320;
 buffer[2426] = 16'h7361;
 buffer[2427] = 16'h2065;
 buffer[2428] = 16'h6F63;
 buffer[2429] = 16'h736E;
 buffer[2430] = 16'h7274;
 buffer[2431] = 16'h6375;
 buffer[2432] = 16'h2E74;
 buffer[2433] = 16'h47C7;
 buffer[2434] = 16'h4963;
 buffer[2435] = 16'h700C;
 buffer[2436] = 16'h12D2;
 buffer[2437] = 16'h24C2;
 buffer[2438] = 16'h0022;
 buffer[2439] = 16'h47C7;
 buffer[2440] = 16'h451E;
 buffer[2441] = 16'h0800;
 buffer[2442] = 16'h130A;
 buffer[2443] = 16'h2EC2;
 buffer[2444] = 16'h0022;
 buffer[2445] = 16'h47C7;
 buffer[2446] = 16'h4528;
 buffer[2447] = 16'h0800;
 buffer[2448] = 16'h1316;
 buffer[2449] = 16'h3E05;
 buffer[2450] = 16'h6F62;
 buffer[2451] = 16'h7964;
 buffer[2452] = 16'h0342;
 buffer[2453] = 16'h1322;
 buffer[2454] = 16'h2844;
 buffer[2455] = 16'h6F74;
 buffer[2456] = 16'h0029;
 buffer[2457] = 16'h6B8D;
 buffer[2458] = 16'h6081;
 buffer[2459] = 16'h4342;
 buffer[2460] = 16'h6147;
 buffer[2461] = 16'h6C00;
 buffer[2462] = 16'h6023;
 buffer[2463] = 16'h710F;
 buffer[2464] = 16'h132C;
 buffer[2465] = 16'h74C2;
 buffer[2466] = 16'h006F;
 buffer[2467] = 16'h47C7;
 buffer[2468] = 16'h4999;
 buffer[2469] = 16'h4787;
 buffer[2470] = 16'h4994;
 buffer[2471] = 16'h0795;
 buffer[2472] = 16'h1342;
 buffer[2473] = 16'h2845;
 buffer[2474] = 16'h742B;
 buffer[2475] = 16'h296F;
 buffer[2476] = 16'h6B8D;
 buffer[2477] = 16'h6081;
 buffer[2478] = 16'h4342;
 buffer[2479] = 16'h6147;
 buffer[2480] = 16'h6C00;
 buffer[2481] = 16'h0367;
 buffer[2482] = 16'h1352;
 buffer[2483] = 16'h2BC3;
 buffer[2484] = 16'h6F74;
 buffer[2485] = 16'h47C7;
 buffer[2486] = 16'h49AC;
 buffer[2487] = 16'h4787;
 buffer[2488] = 16'h4994;
 buffer[2489] = 16'h0795;
 buffer[2490] = 16'h1366;
 buffer[2491] = 16'h670B;
 buffer[2492] = 16'h7465;
 buffer[2493] = 16'h632D;
 buffer[2494] = 16'h7275;
 buffer[2495] = 16'h6572;
 buffer[2496] = 16'h746E;
 buffer[2497] = 16'hFE9A;
 buffer[2498] = 16'h7C0C;
 buffer[2499] = 16'h1376;
 buffer[2500] = 16'h730B;
 buffer[2501] = 16'h7465;
 buffer[2502] = 16'h632D;
 buffer[2503] = 16'h7275;
 buffer[2504] = 16'h6572;
 buffer[2505] = 16'h746E;
 buffer[2506] = 16'hFE9A;
 buffer[2507] = 16'h6023;
 buffer[2508] = 16'h710F;
 buffer[2509] = 16'h1388;
 buffer[2510] = 16'h640B;
 buffer[2511] = 16'h6665;
 buffer[2512] = 16'h6E69;
 buffer[2513] = 16'h7469;
 buffer[2514] = 16'h6F69;
 buffer[2515] = 16'h736E;
 buffer[2516] = 16'hFE90;
 buffer[2517] = 16'h6C00;
 buffer[2518] = 16'h09CA;
 buffer[2519] = 16'h139C;
 buffer[2520] = 16'h3F07;
 buffer[2521] = 16'h6E75;
 buffer[2522] = 16'h7169;
 buffer[2523] = 16'h6575;
 buffer[2524] = 16'h6081;
 buffer[2525] = 16'h49C1;
 buffer[2526] = 16'h4632;
 buffer[2527] = 16'h29E7;
 buffer[2528] = 16'h4528;
 buffer[2529] = 16'h2007;
 buffer[2530] = 16'h6572;
 buffer[2531] = 16'h6564;
 buffer[2532] = 16'h2066;
 buffer[2533] = 16'h6181;
 buffer[2534] = 16'h4523;
 buffer[2535] = 16'h710F;
 buffer[2536] = 16'h13B0;
 buffer[2537] = 16'h3C05;
 buffer[2538] = 16'h2C24;
 buffer[2539] = 16'h3E6E;
 buffer[2540] = 16'h6081;
 buffer[2541] = 16'h417E;
 buffer[2542] = 16'h2A01;
 buffer[2543] = 16'h49DC;
 buffer[2544] = 16'h6081;
 buffer[2545] = 16'h4383;
 buffer[2546] = 16'h6203;
 buffer[2547] = 16'h4392;
 buffer[2548] = 16'hFE9E;
 buffer[2549] = 16'h6023;
 buffer[2550] = 16'h6103;
 buffer[2551] = 16'h6081;
 buffer[2552] = 16'hFEA0;
 buffer[2553] = 16'h6023;
 buffer[2554] = 16'h6103;
 buffer[2555] = 16'h4348;
 buffer[2556] = 16'h49C1;
 buffer[2557] = 16'h6C00;
 buffer[2558] = 16'h6180;
 buffer[2559] = 16'h6023;
 buffer[2560] = 16'h710F;
 buffer[2561] = 16'h6103;
 buffer[2562] = 16'h451E;
 buffer[2563] = 16'h6E04;
 buffer[2564] = 16'h6D61;
 buffer[2565] = 16'h0065;
 buffer[2566] = 16'h06E1;
 buffer[2567] = 16'h13D2;
 buffer[2568] = 16'h2403;
 buffer[2569] = 16'h6E2C;
 buffer[2570] = 16'hFEAC;
 buffer[2571] = 16'h03B3;
 buffer[2572] = 16'h1410;
 buffer[2573] = 16'h2408;
 buffer[2574] = 16'h6F63;
 buffer[2575] = 16'h706D;
 buffer[2576] = 16'h6C69;
 buffer[2577] = 16'h0065;
 buffer[2578] = 16'h4681;
 buffer[2579] = 16'h4277;
 buffer[2580] = 16'h2A1C;
 buffer[2581] = 16'h6C00;
 buffer[2582] = 16'h8080;
 buffer[2583] = 16'h6303;
 buffer[2584] = 16'h2A1B;
 buffer[2585] = 16'h0172;
 buffer[2586] = 16'h0A1C;
 buffer[2587] = 16'h07A1;
 buffer[2588] = 16'h4456;
 buffer[2589] = 16'h2A1F;
 buffer[2590] = 16'h07E7;
 buffer[2591] = 16'h06E1;
 buffer[2592] = 16'h141A;
 buffer[2593] = 16'h6186;
 buffer[2594] = 16'h6F62;
 buffer[2595] = 16'h7472;
 buffer[2596] = 16'h0022;
 buffer[2597] = 16'h47C7;
 buffer[2598] = 16'h46EF;
 buffer[2599] = 16'h0800;
 buffer[2600] = 16'h1442;
 buffer[2601] = 16'h3C07;
 buffer[2602] = 16'h766F;
 buffer[2603] = 16'h7265;
 buffer[2604] = 16'h3E74;
 buffer[2605] = 16'hFEA0;
 buffer[2606] = 16'h6C00;
 buffer[2607] = 16'h49C1;
 buffer[2608] = 16'h6023;
 buffer[2609] = 16'h710F;
 buffer[2610] = 16'h1452;
 buffer[2611] = 16'h6F05;
 buffer[2612] = 16'h6576;
 buffer[2613] = 16'h7472;
 buffer[2614] = 16'hFEAE;
 buffer[2615] = 16'h03B3;
 buffer[2616] = 16'h1466;
 buffer[2617] = 16'h6504;
 buffer[2618] = 16'h6978;
 buffer[2619] = 16'h0074;
 buffer[2620] = 16'h6B8D;
 buffer[2621] = 16'h710F;
 buffer[2622] = 16'h1472;
 buffer[2623] = 16'h3CC3;
 buffer[2624] = 16'h3E3B;
 buffer[2625] = 16'h47C7;
 buffer[2626] = 16'h4A3C;
 buffer[2627] = 16'h4728;
 buffer[2628] = 16'h4A36;
 buffer[2629] = 16'h8000;
 buffer[2630] = 16'h438B;
 buffer[2631] = 16'h6023;
 buffer[2632] = 16'h710F;
 buffer[2633] = 16'h147E;
 buffer[2634] = 16'h3BC1;
 buffer[2635] = 16'hFEB0;
 buffer[2636] = 16'h03B3;
 buffer[2637] = 16'h1494;
 buffer[2638] = 16'h5D01;
 buffer[2639] = 16'h9424;
 buffer[2640] = 16'hFE8A;
 buffer[2641] = 16'h6023;
 buffer[2642] = 16'h710F;
 buffer[2643] = 16'h149C;
 buffer[2644] = 16'h3A01;
 buffer[2645] = 16'h4605;
 buffer[2646] = 16'h4A0A;
 buffer[2647] = 16'h0A4F;
 buffer[2648] = 16'h14A8;
 buffer[2649] = 16'h6909;
 buffer[2650] = 16'h6D6D;
 buffer[2651] = 16'h6465;
 buffer[2652] = 16'h6169;
 buffer[2653] = 16'h6574;
 buffer[2654] = 16'h8080;
 buffer[2655] = 16'hFEA0;
 buffer[2656] = 16'h6C00;
 buffer[2657] = 16'h6C00;
 buffer[2658] = 16'h6403;
 buffer[2659] = 16'hFEA0;
 buffer[2660] = 16'h6C00;
 buffer[2661] = 16'h6023;
 buffer[2662] = 16'h710F;
 buffer[2663] = 16'h14B2;
 buffer[2664] = 16'h7504;
 buffer[2665] = 16'h6573;
 buffer[2666] = 16'h0072;
 buffer[2667] = 16'h4605;
 buffer[2668] = 16'h4A0A;
 buffer[2669] = 16'h4A36;
 buffer[2670] = 16'h47C7;
 buffer[2671] = 16'h41D2;
 buffer[2672] = 16'h0795;
 buffer[2673] = 16'h14D0;
 buffer[2674] = 16'h3C08;
 buffer[2675] = 16'h7263;
 buffer[2676] = 16'h6165;
 buffer[2677] = 16'h6574;
 buffer[2678] = 16'h003E;
 buffer[2679] = 16'h4605;
 buffer[2680] = 16'h4A0A;
 buffer[2681] = 16'h4A36;
 buffer[2682] = 16'h838C;
 buffer[2683] = 16'h07A1;
 buffer[2684] = 16'h14E4;
 buffer[2685] = 16'h6306;
 buffer[2686] = 16'h6572;
 buffer[2687] = 16'h7461;
 buffer[2688] = 16'h0065;
 buffer[2689] = 16'hFEB2;
 buffer[2690] = 16'h03B3;
 buffer[2691] = 16'h14FA;
 buffer[2692] = 16'h7608;
 buffer[2693] = 16'h7261;
 buffer[2694] = 16'h6169;
 buffer[2695] = 16'h6C62;
 buffer[2696] = 16'h0065;
 buffer[2697] = 16'h4A81;
 buffer[2698] = 16'h8000;
 buffer[2699] = 16'h0795;
 buffer[2700] = 16'h1508;
 buffer[2701] = 16'h2847;
 buffer[2702] = 16'h6F64;
 buffer[2703] = 16'h7365;
 buffer[2704] = 16'h293E;
 buffer[2705] = 16'h6B8D;
 buffer[2706] = 16'h8001;
 buffer[2707] = 16'h6903;
 buffer[2708] = 16'h438B;
 buffer[2709] = 16'h8001;
 buffer[2710] = 16'h6903;
 buffer[2711] = 16'hFEA0;
 buffer[2712] = 16'h6C00;
 buffer[2713] = 16'h460B;
 buffer[2714] = 16'h6081;
 buffer[2715] = 16'h4342;
 buffer[2716] = 16'hFFFF;
 buffer[2717] = 16'h6600;
 buffer[2718] = 16'h6403;
 buffer[2719] = 16'h4795;
 buffer[2720] = 16'h6023;
 buffer[2721] = 16'h6103;
 buffer[2722] = 16'h0795;
 buffer[2723] = 16'h151A;
 buffer[2724] = 16'h630C;
 buffer[2725] = 16'h6D6F;
 buffer[2726] = 16'h6970;
 buffer[2727] = 16'h656C;
 buffer[2728] = 16'h6F2D;
 buffer[2729] = 16'h6C6E;
 buffer[2730] = 16'h0079;
 buffer[2731] = 16'h8040;
 buffer[2732] = 16'hFEA0;
 buffer[2733] = 16'h6C00;
 buffer[2734] = 16'h6C00;
 buffer[2735] = 16'h6403;
 buffer[2736] = 16'hFEA0;
 buffer[2737] = 16'h6C00;
 buffer[2738] = 16'h6023;
 buffer[2739] = 16'h710F;
 buffer[2740] = 16'h1548;
 buffer[2741] = 16'h6485;
 buffer[2742] = 16'h656F;
 buffer[2743] = 16'h3E73;
 buffer[2744] = 16'h47C7;
 buffer[2745] = 16'h4A91;
 buffer[2746] = 16'h700C;
 buffer[2747] = 16'h156A;
 buffer[2748] = 16'h6304;
 buffer[2749] = 16'h6168;
 buffer[2750] = 16'h0072;
 buffer[2751] = 16'h4353;
 buffer[2752] = 16'h45FD;
 buffer[2753] = 16'h6310;
 buffer[2754] = 16'h017E;
 buffer[2755] = 16'h1578;
 buffer[2756] = 16'h5B86;
 buffer[2757] = 16'h6863;
 buffer[2758] = 16'h7261;
 buffer[2759] = 16'h005D;
 buffer[2760] = 16'h4ABF;
 buffer[2761] = 16'h07E7;
 buffer[2762] = 16'h1588;
 buffer[2763] = 16'h6308;
 buffer[2764] = 16'h6E6F;
 buffer[2765] = 16'h7473;
 buffer[2766] = 16'h6E61;
 buffer[2767] = 16'h0074;
 buffer[2768] = 16'h4A81;
 buffer[2769] = 16'h4795;
 buffer[2770] = 16'h4A91;
 buffer[2771] = 16'h7C0C;
 buffer[2772] = 16'h1596;
 buffer[2773] = 16'h3209;
 buffer[2774] = 16'h6F63;
 buffer[2775] = 16'h736E;
 buffer[2776] = 16'h6174;
 buffer[2777] = 16'h746E;
 buffer[2778] = 16'h4A81;
 buffer[2779] = 16'h4795;
 buffer[2780] = 16'h4795;
 buffer[2781] = 16'h4AB8;
 buffer[2782] = 16'h037A;
 buffer[2783] = 16'h15AA;
 buffer[2784] = 16'h3209;
 buffer[2785] = 16'h6176;
 buffer[2786] = 16'h6972;
 buffer[2787] = 16'h6261;
 buffer[2788] = 16'h656C;
 buffer[2789] = 16'h4A81;
 buffer[2790] = 16'h8002;
 buffer[2791] = 16'h434E;
 buffer[2792] = 16'h0790;
 buffer[2793] = 16'h15C0;
 buffer[2794] = 16'h6405;
 buffer[2795] = 16'h6665;
 buffer[2796] = 16'h7265;
 buffer[2797] = 16'h4A81;
 buffer[2798] = 16'h8000;
 buffer[2799] = 16'h4795;
 buffer[2800] = 16'h4A91;
 buffer[2801] = 16'h6C00;
 buffer[2802] = 16'h4277;
 buffer[2803] = 16'h8000;
 buffer[2804] = 16'h6703;
 buffer[2805] = 16'h46EF;
 buffer[2806] = 16'h750D;
 buffer[2807] = 16'h696E;
 buffer[2808] = 16'h696E;
 buffer[2809] = 16'h6974;
 buffer[2810] = 16'h6C61;
 buffer[2811] = 16'h7A69;
 buffer[2812] = 16'h6465;
 buffer[2813] = 16'h0172;
 buffer[2814] = 16'h15D4;
 buffer[2815] = 16'h6982;
 buffer[2816] = 16'h0073;
 buffer[2817] = 16'h4787;
 buffer[2818] = 16'h4994;
 buffer[2819] = 16'h6023;
 buffer[2820] = 16'h710F;
 buffer[2821] = 16'h15FE;
 buffer[2822] = 16'h2E03;
 buffer[2823] = 16'h6469;
 buffer[2824] = 16'h4277;
 buffer[2825] = 16'h2B0E;
 buffer[2826] = 16'h4383;
 buffer[2827] = 16'h801F;
 buffer[2828] = 16'h6303;
 buffer[2829] = 16'h04FA;
 buffer[2830] = 16'h450A;
 buffer[2831] = 16'h4528;
 buffer[2832] = 16'h7B08;
 buffer[2833] = 16'h6F6E;
 buffer[2834] = 16'h616E;
 buffer[2835] = 16'h656D;
 buffer[2836] = 16'h007D;
 buffer[2837] = 16'h700C;
 buffer[2838] = 16'h160C;
 buffer[2839] = 16'h7708;
 buffer[2840] = 16'h726F;
 buffer[2841] = 16'h6C64;
 buffer[2842] = 16'h7369;
 buffer[2843] = 16'h0074;
 buffer[2844] = 16'h43A1;
 buffer[2845] = 16'h438B;
 buffer[2846] = 16'h8000;
 buffer[2847] = 16'h4795;
 buffer[2848] = 16'h6081;
 buffer[2849] = 16'hFE9A;
 buffer[2850] = 16'h4342;
 buffer[2851] = 16'h6081;
 buffer[2852] = 16'h6C00;
 buffer[2853] = 16'h4795;
 buffer[2854] = 16'h6023;
 buffer[2855] = 16'h6103;
 buffer[2856] = 16'h8000;
 buffer[2857] = 16'h0795;
 buffer[2858] = 16'h162E;
 buffer[2859] = 16'h6F06;
 buffer[2860] = 16'h6472;
 buffer[2861] = 16'h7265;
 buffer[2862] = 16'h0040;
 buffer[2863] = 16'h6081;
 buffer[2864] = 16'h6C00;
 buffer[2865] = 16'h6081;
 buffer[2866] = 16'h2B39;
 buffer[2867] = 16'h6147;
 buffer[2868] = 16'h4342;
 buffer[2869] = 16'h4B2F;
 buffer[2870] = 16'h6B8D;
 buffer[2871] = 16'h6180;
 buffer[2872] = 16'h731C;
 buffer[2873] = 16'h700F;
 buffer[2874] = 16'h1656;
 buffer[2875] = 16'h6709;
 buffer[2876] = 16'h7465;
 buffer[2877] = 16'h6F2D;
 buffer[2878] = 16'h6472;
 buffer[2879] = 16'h7265;
 buffer[2880] = 16'hFE90;
 buffer[2881] = 16'h0B2F;
 buffer[2882] = 16'h1676;
 buffer[2883] = 16'h3E04;
 buffer[2884] = 16'h6977;
 buffer[2885] = 16'h0064;
 buffer[2886] = 16'h0342;
 buffer[2887] = 16'h1686;
 buffer[2888] = 16'h2E04;
 buffer[2889] = 16'h6977;
 buffer[2890] = 16'h0064;
 buffer[2891] = 16'h44E2;
 buffer[2892] = 16'h6081;
 buffer[2893] = 16'h4B46;
 buffer[2894] = 16'h4342;
 buffer[2895] = 16'h6C00;
 buffer[2896] = 16'h4277;
 buffer[2897] = 16'h2B54;
 buffer[2898] = 16'h4B08;
 buffer[2899] = 16'h710F;
 buffer[2900] = 16'h8000;
 buffer[2901] = 16'h0537;
 buffer[2902] = 16'h1690;
 buffer[2903] = 16'h2104;
 buffer[2904] = 16'h6977;
 buffer[2905] = 16'h0064;
 buffer[2906] = 16'h4B46;
 buffer[2907] = 16'h4342;
 buffer[2908] = 16'hFEA0;
 buffer[2909] = 16'h6C00;
 buffer[2910] = 16'h6180;
 buffer[2911] = 16'h6023;
 buffer[2912] = 16'h710F;
 buffer[2913] = 16'h16AE;
 buffer[2914] = 16'h7604;
 buffer[2915] = 16'h636F;
 buffer[2916] = 16'h0073;
 buffer[2917] = 16'h450A;
 buffer[2918] = 16'h4528;
 buffer[2919] = 16'h7605;
 buffer[2920] = 16'h636F;
 buffer[2921] = 16'h3A73;
 buffer[2922] = 16'hFE9A;
 buffer[2923] = 16'h4342;
 buffer[2924] = 16'h6C00;
 buffer[2925] = 16'h4277;
 buffer[2926] = 16'h2B73;
 buffer[2927] = 16'h6081;
 buffer[2928] = 16'h4B4B;
 buffer[2929] = 16'h4B46;
 buffer[2930] = 16'h0B6C;
 buffer[2931] = 16'h700C;
 buffer[2932] = 16'h16C4;
 buffer[2933] = 16'h6F05;
 buffer[2934] = 16'h6472;
 buffer[2935] = 16'h7265;
 buffer[2936] = 16'h450A;
 buffer[2937] = 16'h4528;
 buffer[2938] = 16'h7307;
 buffer[2939] = 16'h6165;
 buffer[2940] = 16'h6372;
 buffer[2941] = 16'h3A68;
 buffer[2942] = 16'h4B40;
 buffer[2943] = 16'h4277;
 buffer[2944] = 16'h2B85;
 buffer[2945] = 16'h6180;
 buffer[2946] = 16'h4B4B;
 buffer[2947] = 16'h6A00;
 buffer[2948] = 16'h0B7F;
 buffer[2949] = 16'h450A;
 buffer[2950] = 16'h4528;
 buffer[2951] = 16'h6407;
 buffer[2952] = 16'h6665;
 buffer[2953] = 16'h6E69;
 buffer[2954] = 16'h3A65;
 buffer[2955] = 16'h49C1;
 buffer[2956] = 16'h0B4B;
 buffer[2957] = 16'h16EA;
 buffer[2958] = 16'h7309;
 buffer[2959] = 16'h7465;
 buffer[2960] = 16'h6F2D;
 buffer[2961] = 16'h6472;
 buffer[2962] = 16'h7265;
 buffer[2963] = 16'h6081;
 buffer[2964] = 16'h8000;
 buffer[2965] = 16'h6600;
 buffer[2966] = 16'h6703;
 buffer[2967] = 16'h2B9B;
 buffer[2968] = 16'h6103;
 buffer[2969] = 16'hFE94;
 buffer[2970] = 16'h8001;
 buffer[2971] = 16'h8008;
 buffer[2972] = 16'h6181;
 buffer[2973] = 16'h6F03;
 buffer[2974] = 16'h46EF;
 buffer[2975] = 16'h6F12;
 buffer[2976] = 16'h6576;
 buffer[2977] = 16'h2072;
 buffer[2978] = 16'h6973;
 buffer[2979] = 16'h657A;
 buffer[2980] = 16'h6F20;
 buffer[2981] = 16'h2066;
 buffer[2982] = 16'h7623;
 buffer[2983] = 16'h636F;
 buffer[2984] = 16'h0073;
 buffer[2985] = 16'hFE90;
 buffer[2986] = 16'h6180;
 buffer[2987] = 16'h6081;
 buffer[2988] = 16'h2BB6;
 buffer[2989] = 16'h6147;
 buffer[2990] = 16'h6180;
 buffer[2991] = 16'h6181;
 buffer[2992] = 16'h6023;
 buffer[2993] = 16'h6103;
 buffer[2994] = 16'h4342;
 buffer[2995] = 16'h6B8D;
 buffer[2996] = 16'h6A00;
 buffer[2997] = 16'h0BAB;
 buffer[2998] = 16'h6180;
 buffer[2999] = 16'h6023;
 buffer[3000] = 16'h710F;
 buffer[3001] = 16'h171C;
 buffer[3002] = 16'h6F04;
 buffer[3003] = 16'h6C6E;
 buffer[3004] = 16'h0079;
 buffer[3005] = 16'h8000;
 buffer[3006] = 16'h6600;
 buffer[3007] = 16'h0B93;
 buffer[3008] = 16'h1774;
 buffer[3009] = 16'h6104;
 buffer[3010] = 16'h736C;
 buffer[3011] = 16'h006F;
 buffer[3012] = 16'h4B40;
 buffer[3013] = 16'h6181;
 buffer[3014] = 16'h6180;
 buffer[3015] = 16'h6310;
 buffer[3016] = 16'h0B93;
 buffer[3017] = 16'h1782;
 buffer[3018] = 16'h7008;
 buffer[3019] = 16'h6572;
 buffer[3020] = 16'h6976;
 buffer[3021] = 16'h756F;
 buffer[3022] = 16'h0073;
 buffer[3023] = 16'h4B40;
 buffer[3024] = 16'h6180;
 buffer[3025] = 16'h6103;
 buffer[3026] = 16'h6A00;
 buffer[3027] = 16'h0B93;
 buffer[3028] = 16'h1794;
 buffer[3029] = 16'h3E04;
 buffer[3030] = 16'h6F76;
 buffer[3031] = 16'h0063;
 buffer[3032] = 16'h4A81;
 buffer[3033] = 16'h6081;
 buffer[3034] = 16'h4795;
 buffer[3035] = 16'h4B5A;
 buffer[3036] = 16'h4A91;
 buffer[3037] = 16'h6C00;
 buffer[3038] = 16'h6147;
 buffer[3039] = 16'h4B40;
 buffer[3040] = 16'h6180;
 buffer[3041] = 16'h6103;
 buffer[3042] = 16'h6B8D;
 buffer[3043] = 16'h6180;
 buffer[3044] = 16'h0B93;
 buffer[3045] = 16'h17AA;
 buffer[3046] = 16'h7705;
 buffer[3047] = 16'h6469;
 buffer[3048] = 16'h666F;
 buffer[3049] = 16'h4787;
 buffer[3050] = 16'h4994;
 buffer[3051] = 16'h7C0C;
 buffer[3052] = 16'h17CC;
 buffer[3053] = 16'h760A;
 buffer[3054] = 16'h636F;
 buffer[3055] = 16'h6261;
 buffer[3056] = 16'h6C75;
 buffer[3057] = 16'h7261;
 buffer[3058] = 16'h0079;
 buffer[3059] = 16'h4B1C;
 buffer[3060] = 16'h0BD8;
 buffer[3061] = 16'h17DA;
 buffer[3062] = 16'h5F05;
 buffer[3063] = 16'h7974;
 buffer[3064] = 16'h6570;
 buffer[3065] = 16'h6147;
 buffer[3066] = 16'h0BFE;
 buffer[3067] = 16'h4383;
 buffer[3068] = 16'h4359;
 buffer[3069] = 16'h44C8;
 buffer[3070] = 16'h6B81;
 buffer[3071] = 16'h2C04;
 buffer[3072] = 16'h6B8D;
 buffer[3073] = 16'h6A00;
 buffer[3074] = 16'h6147;
 buffer[3075] = 16'h0BFB;
 buffer[3076] = 16'h6B8D;
 buffer[3077] = 16'h6103;
 buffer[3078] = 16'h710F;
 buffer[3079] = 16'h17EC;
 buffer[3080] = 16'h6403;
 buffer[3081] = 16'h2B6D;
 buffer[3082] = 16'h6181;
 buffer[3083] = 16'h8004;
 buffer[3084] = 16'h4537;
 buffer[3085] = 16'h44E2;
 buffer[3086] = 16'h6147;
 buffer[3087] = 16'h0C13;
 buffer[3088] = 16'h4383;
 buffer[3089] = 16'h8003;
 buffer[3090] = 16'h4537;
 buffer[3091] = 16'h6B81;
 buffer[3092] = 16'h2C19;
 buffer[3093] = 16'h6B8D;
 buffer[3094] = 16'h6A00;
 buffer[3095] = 16'h6147;
 buffer[3096] = 16'h0C10;
 buffer[3097] = 16'h6B8D;
 buffer[3098] = 16'h710F;
 buffer[3099] = 16'h1810;
 buffer[3100] = 16'h6404;
 buffer[3101] = 16'h6D75;
 buffer[3102] = 16'h0070;
 buffer[3103] = 16'hFE80;
 buffer[3104] = 16'h6C00;
 buffer[3105] = 16'h6147;
 buffer[3106] = 16'h4429;
 buffer[3107] = 16'h8010;
 buffer[3108] = 16'h430B;
 buffer[3109] = 16'h6147;
 buffer[3110] = 16'h450A;
 buffer[3111] = 16'h8010;
 buffer[3112] = 16'h428C;
 buffer[3113] = 16'h4C0A;
 buffer[3114] = 16'h4156;
 buffer[3115] = 16'h8002;
 buffer[3116] = 16'h44E9;
 buffer[3117] = 16'h4BF9;
 buffer[3118] = 16'h6B81;
 buffer[3119] = 16'h2C34;
 buffer[3120] = 16'h6B8D;
 buffer[3121] = 16'h6A00;
 buffer[3122] = 16'h6147;
 buffer[3123] = 16'h0C26;
 buffer[3124] = 16'h6B8D;
 buffer[3125] = 16'h6103;
 buffer[3126] = 16'h6103;
 buffer[3127] = 16'h6B8D;
 buffer[3128] = 16'hFE80;
 buffer[3129] = 16'h6023;
 buffer[3130] = 16'h710F;
 buffer[3131] = 16'h1838;
 buffer[3132] = 16'h2E02;
 buffer[3133] = 16'h0073;
 buffer[3134] = 16'h450A;
 buffer[3135] = 16'h416A;
 buffer[3136] = 16'h6A00;
 buffer[3137] = 16'h800F;
 buffer[3138] = 16'h6303;
 buffer[3139] = 16'h6147;
 buffer[3140] = 16'h6B81;
 buffer[3141] = 16'h47DB;
 buffer[3142] = 16'h454A;
 buffer[3143] = 16'h6B81;
 buffer[3144] = 16'h2C4D;
 buffer[3145] = 16'h6B8D;
 buffer[3146] = 16'h6A00;
 buffer[3147] = 16'h6147;
 buffer[3148] = 16'h0C44;
 buffer[3149] = 16'h6B8D;
 buffer[3150] = 16'h6103;
 buffer[3151] = 16'h4528;
 buffer[3152] = 16'h3C04;
 buffer[3153] = 16'h6F74;
 buffer[3154] = 16'h0073;
 buffer[3155] = 16'h700C;
 buffer[3156] = 16'h1878;
 buffer[3157] = 16'h2807;
 buffer[3158] = 16'h6E3E;
 buffer[3159] = 16'h6D61;
 buffer[3160] = 16'h2965;
 buffer[3161] = 16'h6C00;
 buffer[3162] = 16'h4277;
 buffer[3163] = 16'h2C63;
 buffer[3164] = 16'h428C;
 buffer[3165] = 16'h460B;
 buffer[3166] = 16'h6503;
 buffer[3167] = 16'h2C62;
 buffer[3168] = 16'h4348;
 buffer[3169] = 16'h0C59;
 buffer[3170] = 16'h700F;
 buffer[3171] = 16'h6103;
 buffer[3172] = 16'h8000;
 buffer[3173] = 16'h700C;
 buffer[3174] = 16'h18AA;
 buffer[3175] = 16'h3E05;
 buffer[3176] = 16'h616E;
 buffer[3177] = 16'h656D;
 buffer[3178] = 16'h6147;
 buffer[3179] = 16'h4B40;
 buffer[3180] = 16'h4277;
 buffer[3181] = 16'h2C86;
 buffer[3182] = 16'h6180;
 buffer[3183] = 16'h6B81;
 buffer[3184] = 16'h6180;
 buffer[3185] = 16'h4C59;
 buffer[3186] = 16'h4277;
 buffer[3187] = 16'h2C84;
 buffer[3188] = 16'h6147;
 buffer[3189] = 16'h6A00;
 buffer[3190] = 16'h6147;
 buffer[3191] = 16'h0C79;
 buffer[3192] = 16'h6103;
 buffer[3193] = 16'h6B81;
 buffer[3194] = 16'h2C7F;
 buffer[3195] = 16'h6B8D;
 buffer[3196] = 16'h6A00;
 buffer[3197] = 16'h6147;
 buffer[3198] = 16'h0C78;
 buffer[3199] = 16'h6B8D;
 buffer[3200] = 16'h6103;
 buffer[3201] = 16'h6B8D;
 buffer[3202] = 16'h6B8D;
 buffer[3203] = 16'h710F;
 buffer[3204] = 16'h6A00;
 buffer[3205] = 16'h0C6C;
 buffer[3206] = 16'h6B8D;
 buffer[3207] = 16'h6103;
 buffer[3208] = 16'h8000;
 buffer[3209] = 16'h700C;
 buffer[3210] = 16'h18CE;
 buffer[3211] = 16'h7303;
 buffer[3212] = 16'h6565;
 buffer[3213] = 16'h4787;
 buffer[3214] = 16'h450A;
 buffer[3215] = 16'h6081;
 buffer[3216] = 16'h6C00;
 buffer[3217] = 16'h4277;
 buffer[3218] = 16'hF00C;
 buffer[3219] = 16'h6503;
 buffer[3220] = 16'h2CA6;
 buffer[3221] = 16'hBFFF;
 buffer[3222] = 16'h6303;
 buffer[3223] = 16'h8001;
 buffer[3224] = 16'h6D03;
 buffer[3225] = 16'h4C6A;
 buffer[3226] = 16'h4277;
 buffer[3227] = 16'h2C9F;
 buffer[3228] = 16'h44E2;
 buffer[3229] = 16'h4B08;
 buffer[3230] = 16'h0CA4;
 buffer[3231] = 16'h6081;
 buffer[3232] = 16'h6C00;
 buffer[3233] = 16'hFFFF;
 buffer[3234] = 16'h6303;
 buffer[3235] = 16'h4543;
 buffer[3236] = 16'h4342;
 buffer[3237] = 16'h0C8F;
 buffer[3238] = 16'h0286;
 buffer[3239] = 16'h1916;
 buffer[3240] = 16'h2807;
 buffer[3241] = 16'h6F77;
 buffer[3242] = 16'h6472;
 buffer[3243] = 16'h2973;
 buffer[3244] = 16'h450A;
 buffer[3245] = 16'h6C00;
 buffer[3246] = 16'h4277;
 buffer[3247] = 16'h2CB5;
 buffer[3248] = 16'h6081;
 buffer[3249] = 16'h4B08;
 buffer[3250] = 16'h44E2;
 buffer[3251] = 16'h4348;
 buffer[3252] = 16'h0CAD;
 buffer[3253] = 16'h700C;
 buffer[3254] = 16'h1950;
 buffer[3255] = 16'h7705;
 buffer[3256] = 16'h726F;
 buffer[3257] = 16'h7364;
 buffer[3258] = 16'h4B40;
 buffer[3259] = 16'h4277;
 buffer[3260] = 16'h2CC8;
 buffer[3261] = 16'h6180;
 buffer[3262] = 16'h450A;
 buffer[3263] = 16'h450A;
 buffer[3264] = 16'h4528;
 buffer[3265] = 16'h3A01;
 buffer[3266] = 16'h6081;
 buffer[3267] = 16'h4B4B;
 buffer[3268] = 16'h450A;
 buffer[3269] = 16'h4CAC;
 buffer[3270] = 16'h6A00;
 buffer[3271] = 16'h0CBB;
 buffer[3272] = 16'h700C;
 buffer[3273] = 16'h196E;
 buffer[3274] = 16'h7603;
 buffer[3275] = 16'h7265;
 buffer[3276] = 16'h8002;
 buffer[3277] = 16'h8100;
 buffer[3278] = 16'h6413;
 buffer[3279] = 16'h8001;
 buffer[3280] = 16'h720F;
 buffer[3281] = 16'h1994;
 buffer[3282] = 16'h6802;
 buffer[3283] = 16'h0069;
 buffer[3284] = 16'h450A;
 buffer[3285] = 16'h4528;
 buffer[3286] = 16'h650B;
 buffer[3287] = 16'h6F66;
 buffer[3288] = 16'h7472;
 buffer[3289] = 16'h2068;
 buffer[3290] = 16'h316A;
 buffer[3291] = 16'h7620;
 buffer[3292] = 16'hFE80;
 buffer[3293] = 16'h6C00;
 buffer[3294] = 16'h4429;
 buffer[3295] = 16'h4CCC;
 buffer[3296] = 16'h43EB;
 buffer[3297] = 16'h43FD;
 buffer[3298] = 16'h43FD;
 buffer[3299] = 16'h802E;
 buffer[3300] = 16'h43F3;
 buffer[3301] = 16'h43FD;
 buffer[3302] = 16'h4415;
 buffer[3303] = 16'h44FA;
 buffer[3304] = 16'hFE80;
 buffer[3305] = 16'h6023;
 buffer[3306] = 16'h6103;
 buffer[3307] = 16'h050A;
 buffer[3308] = 16'h19A4;
 buffer[3309] = 16'h6304;
 buffer[3310] = 16'h6C6F;
 buffer[3311] = 16'h0064;
 buffer[3312] = 16'h8002;
 buffer[3313] = 16'hFE80;
 buffer[3314] = 16'h8042;
 buffer[3315] = 16'h4557;
 buffer[3316] = 16'h476F;
 buffer[3317] = 16'hFE94;
 buffer[3318] = 16'h6081;
 buffer[3319] = 16'hFE90;
 buffer[3320] = 16'h6023;
 buffer[3321] = 16'h6103;
 buffer[3322] = 16'h6081;
 buffer[3323] = 16'hFE9A;
 buffer[3324] = 16'h4370;
 buffer[3325] = 16'h4A36;
 buffer[3326] = 16'hC000;
 buffer[3327] = 16'h4342;
 buffer[3328] = 16'h6081;
 buffer[3329] = 16'h4348;
 buffer[3330] = 16'h6C00;
 buffer[3331] = 16'h4749;
 buffer[3332] = 16'hFEA6;
 buffer[3333] = 16'h43B3;
 buffer[3334] = 16'h4778;
 buffer[3335] = 16'h0CF0;
 buffer[3336] = 16'h19DA;
 buffer[3337] = 16'h3205;
 buffer[3338] = 16'h766F;
 buffer[3339] = 16'h7265;
 buffer[3340] = 16'h6147;
 buffer[3341] = 16'h6147;
 buffer[3342] = 16'h428C;
 buffer[3343] = 16'h6B8D;
 buffer[3344] = 16'h6B8D;
 buffer[3345] = 16'h427E;
 buffer[3346] = 16'h6147;
 buffer[3347] = 16'h427E;
 buffer[3348] = 16'h6B8D;
 buffer[3349] = 16'h700C;
 buffer[3350] = 16'h1A12;
 buffer[3351] = 16'h3205;
 buffer[3352] = 16'h7773;
 buffer[3353] = 16'h7061;
 buffer[3354] = 16'h427E;
 buffer[3355] = 16'h6147;
 buffer[3356] = 16'h427E;
 buffer[3357] = 16'h6B8D;
 buffer[3358] = 16'h700C;
 buffer[3359] = 16'h1A2E;
 buffer[3360] = 16'h3204;
 buffer[3361] = 16'h696E;
 buffer[3362] = 16'h0070;
 buffer[3363] = 16'h427E;
 buffer[3364] = 16'h6103;
 buffer[3365] = 16'h427E;
 buffer[3366] = 16'h710F;
 buffer[3367] = 16'h1A40;
 buffer[3368] = 16'h3204;
 buffer[3369] = 16'h6F72;
 buffer[3370] = 16'h0074;
 buffer[3371] = 16'h6180;
 buffer[3372] = 16'h6147;
 buffer[3373] = 16'h6147;
 buffer[3374] = 16'h4D1A;
 buffer[3375] = 16'h6B8D;
 buffer[3376] = 16'h6B8D;
 buffer[3377] = 16'h6180;
 buffer[3378] = 16'h0D1A;
 buffer[3379] = 16'h1A50;
 buffer[3380] = 16'h6403;
 buffer[3381] = 16'h3D30;
 buffer[3382] = 16'h805F;
 buffer[3383] = 16'h6600;
 buffer[3384] = 16'h4264;
 buffer[3385] = 16'h8043;
 buffer[3386] = 16'h6600;
 buffer[3387] = 16'h7C0C;
 buffer[3388] = 16'h1A68;
 buffer[3389] = 16'h6402;
 buffer[3390] = 16'h003D;
 buffer[3391] = 16'h805F;
 buffer[3392] = 16'h6600;
 buffer[3393] = 16'h4264;
 buffer[3394] = 16'h8041;
 buffer[3395] = 16'h6600;
 buffer[3396] = 16'h7C0C;
 buffer[3397] = 16'h1A7A;
 buffer[3398] = 16'h6402;
 buffer[3399] = 16'h002B;
 buffer[3400] = 16'h805F;
 buffer[3401] = 16'h6600;
 buffer[3402] = 16'h4264;
 buffer[3403] = 16'h805D;
 buffer[3404] = 16'h6600;
 buffer[3405] = 16'h4264;
 buffer[3406] = 16'h805F;
 buffer[3407] = 16'h6600;
 buffer[3408] = 16'h026E;
 buffer[3409] = 16'h1A8C;
 buffer[3410] = 16'h6402;
 buffer[3411] = 16'h002D;
 buffer[3412] = 16'h805D;
 buffer[3413] = 16'h6600;
 buffer[3414] = 16'h4264;
 buffer[3415] = 16'h805F;
 buffer[3416] = 16'h6600;
 buffer[3417] = 16'h4264;
 buffer[3418] = 16'h805D;
 buffer[3419] = 16'h6600;
 buffer[3420] = 16'h026E;
 buffer[3421] = 16'h1AA4;
 buffer[3422] = 16'h7303;
 buffer[3423] = 16'h643E;
 buffer[3424] = 16'h6081;
 buffer[3425] = 16'h791C;
 buffer[3426] = 16'h1ABC;
 buffer[3427] = 16'h6403;
 buffer[3428] = 16'h2B31;
 buffer[3429] = 16'h805F;
 buffer[3430] = 16'h6600;
 buffer[3431] = 16'h4264;
 buffer[3432] = 16'h805B;
 buffer[3433] = 16'h6600;
 buffer[3434] = 16'h026E;
 buffer[3435] = 16'h1AC6;
 buffer[3436] = 16'h6403;
 buffer[3437] = 16'h2D31;
 buffer[3438] = 16'h805F;
 buffer[3439] = 16'h6600;
 buffer[3440] = 16'h4264;
 buffer[3441] = 16'h8059;
 buffer[3442] = 16'h6600;
 buffer[3443] = 16'h026E;
 buffer[3444] = 16'h1AD8;
 buffer[3445] = 16'h6404;
 buffer[3446] = 16'h6F78;
 buffer[3447] = 16'h0072;
 buffer[3448] = 16'h805D;
 buffer[3449] = 16'h6600;
 buffer[3450] = 16'h4264;
 buffer[3451] = 16'h805F;
 buffer[3452] = 16'h6600;
 buffer[3453] = 16'h4264;
 buffer[3454] = 16'h804F;
 buffer[3455] = 16'h6600;
 buffer[3456] = 16'h026E;
 buffer[3457] = 16'h1AEA;
 buffer[3458] = 16'h6404;
 buffer[3459] = 16'h6E61;
 buffer[3460] = 16'h0064;
 buffer[3461] = 16'h805D;
 buffer[3462] = 16'h6600;
 buffer[3463] = 16'h4264;
 buffer[3464] = 16'h805F;
 buffer[3465] = 16'h6600;
 buffer[3466] = 16'h4264;
 buffer[3467] = 16'h804D;
 buffer[3468] = 16'h6600;
 buffer[3469] = 16'h026E;
 buffer[3470] = 16'h1B04;
 buffer[3471] = 16'h6403;
 buffer[3472] = 16'h726F;
 buffer[3473] = 16'h805D;
 buffer[3474] = 16'h6600;
 buffer[3475] = 16'h4264;
 buffer[3476] = 16'h805F;
 buffer[3477] = 16'h6600;
 buffer[3478] = 16'h4264;
 buffer[3479] = 16'h804B;
 buffer[3480] = 16'h6600;
 buffer[3481] = 16'h026E;
 buffer[3482] = 16'h1B1E;
 buffer[3483] = 16'h6407;
 buffer[3484] = 16'h6E69;
 buffer[3485] = 16'h6576;
 buffer[3486] = 16'h7472;
 buffer[3487] = 16'h805F;
 buffer[3488] = 16'h6600;
 buffer[3489] = 16'h4264;
 buffer[3490] = 16'h8051;
 buffer[3491] = 16'h6600;
 buffer[3492] = 16'h026E;
 buffer[3493] = 16'h1B36;
 buffer[3494] = 16'h6403;
 buffer[3495] = 16'h2A32;
 buffer[3496] = 16'h805F;
 buffer[3497] = 16'h6600;
 buffer[3498] = 16'h4264;
 buffer[3499] = 16'h8057;
 buffer[3500] = 16'h6600;
 buffer[3501] = 16'h026E;
 buffer[3502] = 16'h1B4C;
 buffer[3503] = 16'h6403;
 buffer[3504] = 16'h2F32;
 buffer[3505] = 16'h805F;
 buffer[3506] = 16'h6600;
 buffer[3507] = 16'h4264;
 buffer[3508] = 16'h8055;
 buffer[3509] = 16'h6600;
 buffer[3510] = 16'h026E;
 buffer[3511] = 16'h1B5E;
 buffer[3512] = 16'h6404;
 buffer[3513] = 16'h6261;
 buffer[3514] = 16'h0073;
 buffer[3515] = 16'h805F;
 buffer[3516] = 16'h6600;
 buffer[3517] = 16'h4264;
 buffer[3518] = 16'h8049;
 buffer[3519] = 16'h6600;
 buffer[3520] = 16'h026E;
 buffer[3521] = 16'h1B70;
 buffer[3522] = 16'h6404;
 buffer[3523] = 16'h616D;
 buffer[3524] = 16'h0078;
 buffer[3525] = 16'h805D;
 buffer[3526] = 16'h6600;
 buffer[3527] = 16'h4264;
 buffer[3528] = 16'h805F;
 buffer[3529] = 16'h6600;
 buffer[3530] = 16'h4264;
 buffer[3531] = 16'h8047;
 buffer[3532] = 16'h6600;
 buffer[3533] = 16'h026E;
 buffer[3534] = 16'h1B84;
 buffer[3535] = 16'h6404;
 buffer[3536] = 16'h696D;
 buffer[3537] = 16'h006E;
 buffer[3538] = 16'h805D;
 buffer[3539] = 16'h6600;
 buffer[3540] = 16'h4264;
 buffer[3541] = 16'h805F;
 buffer[3542] = 16'h6600;
 buffer[3543] = 16'h4264;
 buffer[3544] = 16'h8045;
 buffer[3545] = 16'h6600;
 buffer[3546] = 16'h026E;
 buffer[3547] = 16'h1B9E;
 buffer[3548] = 16'h6C04;
 buffer[3549] = 16'h6465;
 buffer[3550] = 16'h0040;
 buffer[3551] = 16'h8FFD;
 buffer[3552] = 16'h6600;
 buffer[3553] = 16'h7C0C;
 buffer[3554] = 16'h1BB8;
 buffer[3555] = 16'h6C04;
 buffer[3556] = 16'h6465;
 buffer[3557] = 16'h0021;
 buffer[3558] = 16'h8FFD;
 buffer[3559] = 16'h6600;
 buffer[3560] = 16'h6023;
 buffer[3561] = 16'h710F;
 buffer[3562] = 16'h1BC6;
 buffer[3563] = 16'h6208;
 buffer[3564] = 16'h7475;
 buffer[3565] = 16'h6F74;
 buffer[3566] = 16'h736E;
 buffer[3567] = 16'h0040;
 buffer[3568] = 16'h8FFC;
 buffer[3569] = 16'h6600;
 buffer[3570] = 16'h7C0C;
 buffer[3571] = 16'h1BD6;
 buffer[3572] = 16'h6205;
 buffer[3573] = 16'h6565;
 buffer[3574] = 16'h2170;
 buffer[3575] = 16'h6081;
 buffer[3576] = 16'h801D;
 buffer[3577] = 16'h6600;
 buffer[3578] = 16'h6023;
 buffer[3579] = 16'h6103;
 buffer[3580] = 16'h8019;
 buffer[3581] = 16'h6600;
 buffer[3582] = 16'h6023;
 buffer[3583] = 16'h6103;
 buffer[3584] = 16'h6081;
 buffer[3585] = 16'h801E;
 buffer[3586] = 16'h6600;
 buffer[3587] = 16'h6023;
 buffer[3588] = 16'h6103;
 buffer[3589] = 16'h801A;
 buffer[3590] = 16'h6600;
 buffer[3591] = 16'h6023;
 buffer[3592] = 16'h6103;
 buffer[3593] = 16'h6081;
 buffer[3594] = 16'h801F;
 buffer[3595] = 16'h6600;
 buffer[3596] = 16'h6023;
 buffer[3597] = 16'h6103;
 buffer[3598] = 16'h801B;
 buffer[3599] = 16'h6600;
 buffer[3600] = 16'h6023;
 buffer[3601] = 16'h6103;
 buffer[3602] = 16'h6081;
 buffer[3603] = 16'h801C;
 buffer[3604] = 16'h6600;
 buffer[3605] = 16'h6023;
 buffer[3606] = 16'h6103;
 buffer[3607] = 16'h8018;
 buffer[3608] = 16'h6600;
 buffer[3609] = 16'h6023;
 buffer[3610] = 16'h710F;
 buffer[3611] = 16'h1BE8;
 buffer[3612] = 16'h6205;
 buffer[3613] = 16'h6565;
 buffer[3614] = 16'h3F70;
 buffer[3615] = 16'h801C;
 buffer[3616] = 16'h6600;
 buffer[3617] = 16'h6C00;
 buffer[3618] = 16'h6010;
 buffer[3619] = 16'h2E1F;
 buffer[3620] = 16'h8018;
 buffer[3621] = 16'h6600;
 buffer[3622] = 16'h6C00;
 buffer[3623] = 16'h6010;
 buffer[3624] = 16'h2E24;
 buffer[3625] = 16'h700C;
 buffer[3626] = 16'h1C38;
 buffer[3627] = 16'h6206;
 buffer[3628] = 16'h6565;
 buffer[3629] = 16'h4C70;
 buffer[3630] = 16'h0021;
 buffer[3631] = 16'h801D;
 buffer[3632] = 16'h6600;
 buffer[3633] = 16'h6023;
 buffer[3634] = 16'h6103;
 buffer[3635] = 16'h801E;
 buffer[3636] = 16'h6600;
 buffer[3637] = 16'h6023;
 buffer[3638] = 16'h6103;
 buffer[3639] = 16'h801F;
 buffer[3640] = 16'h6600;
 buffer[3641] = 16'h6023;
 buffer[3642] = 16'h6103;
 buffer[3643] = 16'h801C;
 buffer[3644] = 16'h6600;
 buffer[3645] = 16'h6023;
 buffer[3646] = 16'h710F;
 buffer[3647] = 16'h1C56;
 buffer[3648] = 16'h6206;
 buffer[3649] = 16'h6565;
 buffer[3650] = 16'h5270;
 buffer[3651] = 16'h0021;
 buffer[3652] = 16'h8019;
 buffer[3653] = 16'h6600;
 buffer[3654] = 16'h6023;
 buffer[3655] = 16'h6103;
 buffer[3656] = 16'h801A;
 buffer[3657] = 16'h6600;
 buffer[3658] = 16'h6023;
 buffer[3659] = 16'h6103;
 buffer[3660] = 16'h801B;
 buffer[3661] = 16'h6600;
 buffer[3662] = 16'h6023;
 buffer[3663] = 16'h6103;
 buffer[3664] = 16'h8018;
 buffer[3665] = 16'h6600;
 buffer[3666] = 16'h6023;
 buffer[3667] = 16'h710F;
 buffer[3668] = 16'h1C80;
 buffer[3669] = 16'h6206;
 buffer[3670] = 16'h6565;
 buffer[3671] = 16'h4C70;
 buffer[3672] = 16'h003F;
 buffer[3673] = 16'h801C;
 buffer[3674] = 16'h6600;
 buffer[3675] = 16'h6C00;
 buffer[3676] = 16'h6010;
 buffer[3677] = 16'h2E59;
 buffer[3678] = 16'h700C;
 buffer[3679] = 16'h1CAA;
 buffer[3680] = 16'h6206;
 buffer[3681] = 16'h6565;
 buffer[3682] = 16'h5270;
 buffer[3683] = 16'h003F;
 buffer[3684] = 16'h8018;
 buffer[3685] = 16'h6600;
 buffer[3686] = 16'h6C00;
 buffer[3687] = 16'h6010;
 buffer[3688] = 16'h2E64;
 buffer[3689] = 16'h700C;
 buffer[3690] = 16'h1CC0;
 buffer[3691] = 16'h6306;
 buffer[3692] = 16'h6F6C;
 buffer[3693] = 16'h6B63;
 buffer[3694] = 16'h0040;
 buffer[3695] = 16'h8FFB;
 buffer[3696] = 16'h6600;
 buffer[3697] = 16'h7C0C;
 buffer[3698] = 16'h1CD6;
 buffer[3699] = 16'h7409;
 buffer[3700] = 16'h6D69;
 buffer[3701] = 16'h7265;
 buffer[3702] = 16'h6831;
 buffer[3703] = 16'h217A;
 buffer[3704] = 16'h8001;
 buffer[3705] = 16'h8012;
 buffer[3706] = 16'h6600;
 buffer[3707] = 16'h6023;
 buffer[3708] = 16'h710F;
 buffer[3709] = 16'h1CE6;
 buffer[3710] = 16'h7409;
 buffer[3711] = 16'h6D69;
 buffer[3712] = 16'h7265;
 buffer[3713] = 16'h6831;
 buffer[3714] = 16'h407A;
 buffer[3715] = 16'h8012;
 buffer[3716] = 16'h6600;
 buffer[3717] = 16'h7C0C;
 buffer[3718] = 16'h1CFC;
 buffer[3719] = 16'h740A;
 buffer[3720] = 16'h6D69;
 buffer[3721] = 16'h7265;
 buffer[3722] = 16'h6B31;
 buffer[3723] = 16'h7A68;
 buffer[3724] = 16'h0021;
 buffer[3725] = 16'h8011;
 buffer[3726] = 16'h6600;
 buffer[3727] = 16'h6023;
 buffer[3728] = 16'h710F;
 buffer[3729] = 16'h1D0E;
 buffer[3730] = 16'h740A;
 buffer[3731] = 16'h6D69;
 buffer[3732] = 16'h7265;
 buffer[3733] = 16'h6B31;
 buffer[3734] = 16'h7A68;
 buffer[3735] = 16'h0040;
 buffer[3736] = 16'h8011;
 buffer[3737] = 16'h6600;
 buffer[3738] = 16'h7C0C;
 buffer[3739] = 16'h1D24;
 buffer[3740] = 16'h740A;
 buffer[3741] = 16'h6D69;
 buffer[3742] = 16'h7265;
 buffer[3743] = 16'h6B31;
 buffer[3744] = 16'h7A68;
 buffer[3745] = 16'h003F;
 buffer[3746] = 16'h8011;
 buffer[3747] = 16'h6600;
 buffer[3748] = 16'h6C00;
 buffer[3749] = 16'h6010;
 buffer[3750] = 16'h2EA2;
 buffer[3751] = 16'h700C;
 buffer[3752] = 16'h1D38;
 buffer[3753] = 16'h7305;
 buffer[3754] = 16'h656C;
 buffer[3755] = 16'h7065;
 buffer[3756] = 16'h8010;
 buffer[3757] = 16'h6600;
 buffer[3758] = 16'h6023;
 buffer[3759] = 16'h6103;
 buffer[3760] = 16'h8010;
 buffer[3761] = 16'h6600;
 buffer[3762] = 16'h6C00;
 buffer[3763] = 16'h6010;
 buffer[3764] = 16'h2EB0;
 buffer[3765] = 16'h700C;
 buffer[3766] = 16'h1D52;
 buffer[3767] = 16'h7203;
 buffer[3768] = 16'h676E;
 buffer[3769] = 16'h801F;
 buffer[3770] = 16'h6600;
 buffer[3771] = 16'h6C00;
 buffer[3772] = 16'h6180;
 buffer[3773] = 16'h42F8;
 buffer[3774] = 16'h710F;
 buffer[3775] = 16'h1D6E;
 buffer[3776] = 16'h7607;
 buffer[3777] = 16'h6C62;
 buffer[3778] = 16'h6E61;
 buffer[3779] = 16'h3F6B;
 buffer[3780] = 16'h8000;
 buffer[3781] = 16'h6600;
 buffer[3782] = 16'h6C00;
 buffer[3783] = 16'h6110;
 buffer[3784] = 16'h2EC4;
 buffer[3785] = 16'h700C;
 buffer[3786] = 16'h1D80;
 buffer[3787] = 16'h620B;
 buffer[3788] = 16'h6361;
 buffer[3789] = 16'h676B;
 buffer[3790] = 16'h6F72;
 buffer[3791] = 16'h6E75;
 buffer[3792] = 16'h2164;
 buffer[3793] = 16'h800D;
 buffer[3794] = 16'h6600;
 buffer[3795] = 16'h6023;
 buffer[3796] = 16'h6103;
 buffer[3797] = 16'h800E;
 buffer[3798] = 16'h6600;
 buffer[3799] = 16'h6023;
 buffer[3800] = 16'h6103;
 buffer[3801] = 16'h800F;
 buffer[3802] = 16'h6600;
 buffer[3803] = 16'h6023;
 buffer[3804] = 16'h710F;
 buffer[3805] = 16'h1D96;
 buffer[3806] = 16'h6704;
 buffer[3807] = 16'h7570;
 buffer[3808] = 16'h003F;
 buffer[3809] = 16'h80F8;
 buffer[3810] = 16'h6600;
 buffer[3811] = 16'h6C00;
 buffer[3812] = 16'h6010;
 buffer[3813] = 16'h2EE1;
 buffer[3814] = 16'h700C;
 buffer[3815] = 16'h1DBC;
 buffer[3816] = 16'h6704;
 buffer[3817] = 16'h7570;
 buffer[3818] = 16'h0021;
 buffer[3819] = 16'h4EE1;
 buffer[3820] = 16'h80F8;
 buffer[3821] = 16'h6600;
 buffer[3822] = 16'h6023;
 buffer[3823] = 16'h710F;
 buffer[3824] = 16'h1DD0;
 buffer[3825] = 16'h7006;
 buffer[3826] = 16'h7869;
 buffer[3827] = 16'h6C65;
 buffer[3828] = 16'h0021;
 buffer[3829] = 16'h80FE;
 buffer[3830] = 16'h6600;
 buffer[3831] = 16'h6023;
 buffer[3832] = 16'h6103;
 buffer[3833] = 16'h80FF;
 buffer[3834] = 16'h6600;
 buffer[3835] = 16'h6023;
 buffer[3836] = 16'h6103;
 buffer[3837] = 16'h80FD;
 buffer[3838] = 16'h6600;
 buffer[3839] = 16'h6023;
 buffer[3840] = 16'h6103;
 buffer[3841] = 16'h8001;
 buffer[3842] = 16'h0EEB;
 buffer[3843] = 16'h1DE2;
 buffer[3844] = 16'h720A;
 buffer[3845] = 16'h6365;
 buffer[3846] = 16'h6174;
 buffer[3847] = 16'h676E;
 buffer[3848] = 16'h656C;
 buffer[3849] = 16'h0021;
 buffer[3850] = 16'h80FB;
 buffer[3851] = 16'h6600;
 buffer[3852] = 16'h6023;
 buffer[3853] = 16'h6103;
 buffer[3854] = 16'h80FC;
 buffer[3855] = 16'h6600;
 buffer[3856] = 16'h6023;
 buffer[3857] = 16'h6103;
 buffer[3858] = 16'h80FE;
 buffer[3859] = 16'h6600;
 buffer[3860] = 16'h6023;
 buffer[3861] = 16'h6103;
 buffer[3862] = 16'h80FF;
 buffer[3863] = 16'h6600;
 buffer[3864] = 16'h6023;
 buffer[3865] = 16'h6103;
 buffer[3866] = 16'h80FD;
 buffer[3867] = 16'h6600;
 buffer[3868] = 16'h6023;
 buffer[3869] = 16'h6103;
 buffer[3870] = 16'h8002;
 buffer[3871] = 16'h0EEB;
 buffer[3872] = 16'h1E08;
 buffer[3873] = 16'h6C05;
 buffer[3874] = 16'h6E69;
 buffer[3875] = 16'h2165;
 buffer[3876] = 16'h80FB;
 buffer[3877] = 16'h6600;
 buffer[3878] = 16'h6023;
 buffer[3879] = 16'h6103;
 buffer[3880] = 16'h80FC;
 buffer[3881] = 16'h6600;
 buffer[3882] = 16'h6023;
 buffer[3883] = 16'h6103;
 buffer[3884] = 16'h80FE;
 buffer[3885] = 16'h6600;
 buffer[3886] = 16'h6023;
 buffer[3887] = 16'h6103;
 buffer[3888] = 16'h80FF;
 buffer[3889] = 16'h6600;
 buffer[3890] = 16'h6023;
 buffer[3891] = 16'h6103;
 buffer[3892] = 16'h80FD;
 buffer[3893] = 16'h6600;
 buffer[3894] = 16'h6023;
 buffer[3895] = 16'h6103;
 buffer[3896] = 16'h8003;
 buffer[3897] = 16'h0EEB;
 buffer[3898] = 16'h1E42;
 buffer[3899] = 16'h6307;
 buffer[3900] = 16'h7269;
 buffer[3901] = 16'h6C63;
 buffer[3902] = 16'h2165;
 buffer[3903] = 16'h80FC;
 buffer[3904] = 16'h6600;
 buffer[3905] = 16'h6023;
 buffer[3906] = 16'h6103;
 buffer[3907] = 16'h80FE;
 buffer[3908] = 16'h6600;
 buffer[3909] = 16'h6023;
 buffer[3910] = 16'h6103;
 buffer[3911] = 16'h80FF;
 buffer[3912] = 16'h6600;
 buffer[3913] = 16'h6023;
 buffer[3914] = 16'h6103;
 buffer[3915] = 16'h80FD;
 buffer[3916] = 16'h6600;
 buffer[3917] = 16'h6023;
 buffer[3918] = 16'h6103;
 buffer[3919] = 16'h8004;
 buffer[3920] = 16'h0EEB;
 buffer[3921] = 16'h1E76;
 buffer[3922] = 16'h6608;
 buffer[3923] = 16'h6963;
 buffer[3924] = 16'h6372;
 buffer[3925] = 16'h656C;
 buffer[3926] = 16'h0021;
 buffer[3927] = 16'h80FC;
 buffer[3928] = 16'h6600;
 buffer[3929] = 16'h6023;
 buffer[3930] = 16'h6103;
 buffer[3931] = 16'h80FE;
 buffer[3932] = 16'h6600;
 buffer[3933] = 16'h6023;
 buffer[3934] = 16'h6103;
 buffer[3935] = 16'h80FF;
 buffer[3936] = 16'h6600;
 buffer[3937] = 16'h6023;
 buffer[3938] = 16'h6103;
 buffer[3939] = 16'h80FD;
 buffer[3940] = 16'h6600;
 buffer[3941] = 16'h6023;
 buffer[3942] = 16'h6103;
 buffer[3943] = 16'h8006;
 buffer[3944] = 16'h0EEB;
 buffer[3945] = 16'h1EA4;
 buffer[3946] = 16'h7409;
 buffer[3947] = 16'h6972;
 buffer[3948] = 16'h6E61;
 buffer[3949] = 16'h6C67;
 buffer[3950] = 16'h2165;
 buffer[3951] = 16'h80F9;
 buffer[3952] = 16'h6600;
 buffer[3953] = 16'h6023;
 buffer[3954] = 16'h6103;
 buffer[3955] = 16'h80FA;
 buffer[3956] = 16'h6600;
 buffer[3957] = 16'h6023;
 buffer[3958] = 16'h6103;
 buffer[3959] = 16'h80FB;
 buffer[3960] = 16'h6600;
 buffer[3961] = 16'h6023;
 buffer[3962] = 16'h6103;
 buffer[3963] = 16'h80FC;
 buffer[3964] = 16'h6600;
 buffer[3965] = 16'h6023;
 buffer[3966] = 16'h6103;
 buffer[3967] = 16'h80FE;
 buffer[3968] = 16'h6600;
 buffer[3969] = 16'h6023;
 buffer[3970] = 16'h6103;
 buffer[3971] = 16'h80FF;
 buffer[3972] = 16'h6600;
 buffer[3973] = 16'h6023;
 buffer[3974] = 16'h6103;
 buffer[3975] = 16'h80FD;
 buffer[3976] = 16'h6600;
 buffer[3977] = 16'h6023;
 buffer[3978] = 16'h6103;
 buffer[3979] = 16'h8007;
 buffer[3980] = 16'h0EEB;
 buffer[3981] = 16'h1ED4;
 buffer[3982] = 16'h6206;
 buffer[3983] = 16'h696C;
 buffer[3984] = 16'h3174;
 buffer[3985] = 16'h0021;
 buffer[3986] = 16'h80FE;
 buffer[3987] = 16'h6600;
 buffer[3988] = 16'h6023;
 buffer[3989] = 16'h6103;
 buffer[3990] = 16'h80FF;
 buffer[3991] = 16'h6600;
 buffer[3992] = 16'h6023;
 buffer[3993] = 16'h6103;
 buffer[3994] = 16'h80FC;
 buffer[3995] = 16'h6600;
 buffer[3996] = 16'h6023;
 buffer[3997] = 16'h6103;
 buffer[3998] = 16'h80FD;
 buffer[3999] = 16'h6600;
 buffer[4000] = 16'h6023;
 buffer[4001] = 16'h6103;
 buffer[4002] = 16'h8005;
 buffer[4003] = 16'h0EEB;
 buffer[4004] = 16'h1F1C;
 buffer[4005] = 16'h620A;
 buffer[4006] = 16'h696C;
 buffer[4007] = 16'h3174;
 buffer[4008] = 16'h6974;
 buffer[4009] = 16'h656C;
 buffer[4010] = 16'h0021;
 buffer[4011] = 16'h80F4;
 buffer[4012] = 16'h6600;
 buffer[4013] = 16'h6023;
 buffer[4014] = 16'h6103;
 buffer[4015] = 16'h8010;
 buffer[4016] = 16'h6A00;
 buffer[4017] = 16'h6081;
 buffer[4018] = 16'h80F3;
 buffer[4019] = 16'h6600;
 buffer[4020] = 16'h6023;
 buffer[4021] = 16'h6103;
 buffer[4022] = 16'h6180;
 buffer[4023] = 16'h80F2;
 buffer[4024] = 16'h6600;
 buffer[4025] = 16'h6023;
 buffer[4026] = 16'h6103;
 buffer[4027] = 16'h6081;
 buffer[4028] = 16'h6010;
 buffer[4029] = 16'h2FB0;
 buffer[4030] = 16'h710F;
 buffer[4031] = 16'h1F4A;
 buffer[4032] = 16'h6303;
 buffer[4033] = 16'h2173;
 buffer[4034] = 16'h8005;
 buffer[4035] = 16'h80F7;
 buffer[4036] = 16'h6600;
 buffer[4037] = 16'h6023;
 buffer[4038] = 16'h6103;
 buffer[4039] = 16'h8040;
 buffer[4040] = 16'h8000;
 buffer[4041] = 16'h8000;
 buffer[4042] = 16'h82F7;
 buffer[4043] = 16'h81DF;
 buffer[4044] = 16'h0F0A;
 buffer[4045] = 16'h1F80;
 buffer[4046] = 16'h6C08;
 buffer[4047] = 16'h6C73;
 buffer[4048] = 16'h6974;
 buffer[4049] = 16'h656C;
 buffer[4050] = 16'h0021;
 buffer[4051] = 16'h80C7;
 buffer[4052] = 16'h6600;
 buffer[4053] = 16'h6023;
 buffer[4054] = 16'h6103;
 buffer[4055] = 16'h8080;
 buffer[4056] = 16'h6A00;
 buffer[4057] = 16'h6081;
 buffer[4058] = 16'h80C6;
 buffer[4059] = 16'h6600;
 buffer[4060] = 16'h6023;
 buffer[4061] = 16'h6103;
 buffer[4062] = 16'h6180;
 buffer[4063] = 16'h80C5;
 buffer[4064] = 16'h6600;
 buffer[4065] = 16'h6023;
 buffer[4066] = 16'h6103;
 buffer[4067] = 16'h6081;
 buffer[4068] = 16'h6010;
 buffer[4069] = 16'h2FD8;
 buffer[4070] = 16'h710F;
 buffer[4071] = 16'h1F9C;
 buffer[4072] = 16'h6C0A;
 buffer[4073] = 16'h6C73;
 buffer[4074] = 16'h7073;
 buffer[4075] = 16'h6972;
 buffer[4076] = 16'h6574;
 buffer[4077] = 16'h0021;
 buffer[4078] = 16'h80CF;
 buffer[4079] = 16'h6600;
 buffer[4080] = 16'h6023;
 buffer[4081] = 16'h6103;
 buffer[4082] = 16'h80C9;
 buffer[4083] = 16'h6600;
 buffer[4084] = 16'h6023;
 buffer[4085] = 16'h6103;
 buffer[4086] = 16'h80CE;
 buffer[4087] = 16'h6600;
 buffer[4088] = 16'h6023;
 buffer[4089] = 16'h6103;
 buffer[4090] = 16'h80CD;
 buffer[4091] = 16'h6600;
 buffer[4092] = 16'h6023;
 buffer[4093] = 16'h6103;
 buffer[4094] = 16'h80CA;
 buffer[4095] = 16'h6600;
 buffer[4096] = 16'h6023;
 buffer[4097] = 16'h6103;
 buffer[4098] = 16'h80CB;
 buffer[4099] = 16'h6600;
 buffer[4100] = 16'h6023;
 buffer[4101] = 16'h6103;
 buffer[4102] = 16'h80CC;
 buffer[4103] = 16'h6600;
 buffer[4104] = 16'h6023;
 buffer[4105] = 16'h710F;
 buffer[4106] = 16'h1FD0;
 buffer[4107] = 16'h6C0A;
 buffer[4108] = 16'h6C73;
 buffer[4109] = 16'h7075;
 buffer[4110] = 16'h6164;
 buffer[4111] = 16'h6574;
 buffer[4112] = 16'h0021;
 buffer[4113] = 16'h80CF;
 buffer[4114] = 16'h6600;
 buffer[4115] = 16'h6023;
 buffer[4116] = 16'h6103;
 buffer[4117] = 16'h80C1;
 buffer[4118] = 16'h6600;
 buffer[4119] = 16'h6023;
 buffer[4120] = 16'h710F;
 buffer[4121] = 16'h2016;
 buffer[4122] = 16'h7508;
 buffer[4123] = 16'h6C73;
 buffer[4124] = 16'h6974;
 buffer[4125] = 16'h656C;
 buffer[4126] = 16'h0021;
 buffer[4127] = 16'h80B7;
 buffer[4128] = 16'h6600;
 buffer[4129] = 16'h6023;
 buffer[4130] = 16'h6103;
 buffer[4131] = 16'h8080;
 buffer[4132] = 16'h6A00;
 buffer[4133] = 16'h6081;
 buffer[4134] = 16'h80B6;
 buffer[4135] = 16'h6600;
 buffer[4136] = 16'h6023;
 buffer[4137] = 16'h6103;
 buffer[4138] = 16'h6180;
 buffer[4139] = 16'h80B5;
 buffer[4140] = 16'h6600;
 buffer[4141] = 16'h6023;
 buffer[4142] = 16'h6103;
 buffer[4143] = 16'h6081;
 buffer[4144] = 16'h6010;
 buffer[4145] = 16'h3024;
 buffer[4146] = 16'h710F;
 buffer[4147] = 16'h2034;
 buffer[4148] = 16'h750A;
 buffer[4149] = 16'h6C73;
 buffer[4150] = 16'h7073;
 buffer[4151] = 16'h6972;
 buffer[4152] = 16'h6574;
 buffer[4153] = 16'h0021;
 buffer[4154] = 16'h80BF;
 buffer[4155] = 16'h6600;
 buffer[4156] = 16'h6023;
 buffer[4157] = 16'h6103;
 buffer[4158] = 16'h80B9;
 buffer[4159] = 16'h6600;
 buffer[4160] = 16'h6023;
 buffer[4161] = 16'h6103;
 buffer[4162] = 16'h80BE;
 buffer[4163] = 16'h6600;
 buffer[4164] = 16'h6023;
 buffer[4165] = 16'h6103;
 buffer[4166] = 16'h80BD;
 buffer[4167] = 16'h6600;
 buffer[4168] = 16'h6023;
 buffer[4169] = 16'h6103;
 buffer[4170] = 16'h80BA;
 buffer[4171] = 16'h6600;
 buffer[4172] = 16'h6023;
 buffer[4173] = 16'h6103;
 buffer[4174] = 16'h80BB;
 buffer[4175] = 16'h6600;
 buffer[4176] = 16'h6023;
 buffer[4177] = 16'h6103;
 buffer[4178] = 16'h80BC;
 buffer[4179] = 16'h6600;
 buffer[4180] = 16'h6023;
 buffer[4181] = 16'h710F;
 buffer[4182] = 16'h2068;
 buffer[4183] = 16'h750A;
 buffer[4184] = 16'h6C73;
 buffer[4185] = 16'h7075;
 buffer[4186] = 16'h6164;
 buffer[4187] = 16'h6574;
 buffer[4188] = 16'h0021;
 buffer[4189] = 16'h80BF;
 buffer[4190] = 16'h6600;
 buffer[4191] = 16'h6023;
 buffer[4192] = 16'h6103;
 buffer[4193] = 16'h80B1;
 buffer[4194] = 16'h6600;
 buffer[4195] = 16'h6023;
 buffer[4196] = 16'h710F;
 buffer[4197] = 16'h20AE;
 buffer[4198] = 16'h760D;
 buffer[4199] = 16'h6365;
 buffer[4200] = 16'h6F74;
 buffer[4201] = 16'h7672;
 buffer[4202] = 16'h7265;
 buffer[4203] = 16'h6574;
 buffer[4204] = 16'h2178;
 buffer[4205] = 16'h8089;
 buffer[4206] = 16'h6600;
 buffer[4207] = 16'h6023;
 buffer[4208] = 16'h6103;
 buffer[4209] = 16'h808A;
 buffer[4210] = 16'h6600;
 buffer[4211] = 16'h6023;
 buffer[4212] = 16'h6103;
 buffer[4213] = 16'h8087;
 buffer[4214] = 16'h6600;
 buffer[4215] = 16'h6023;
 buffer[4216] = 16'h6103;
 buffer[4217] = 16'h8088;
 buffer[4218] = 16'h6600;
 buffer[4219] = 16'h6023;
 buffer[4220] = 16'h6103;
 buffer[4221] = 16'h8086;
 buffer[4222] = 16'h6600;
 buffer[4223] = 16'h6023;
 buffer[4224] = 16'h710F;
 buffer[4225] = 16'h20CC;
 buffer[4226] = 16'h7607;
 buffer[4227] = 16'h6365;
 buffer[4228] = 16'h6F74;
 buffer[4229] = 16'h3F72;
 buffer[4230] = 16'h808B;
 buffer[4231] = 16'h6600;
 buffer[4232] = 16'h6C00;
 buffer[4233] = 16'h6010;
 buffer[4234] = 16'h3086;
 buffer[4235] = 16'h700C;
 buffer[4236] = 16'h2104;
 buffer[4237] = 16'h7607;
 buffer[4238] = 16'h6365;
 buffer[4239] = 16'h6F74;
 buffer[4240] = 16'h2172;
 buffer[4241] = 16'h5086;
 buffer[4242] = 16'h808F;
 buffer[4243] = 16'h6600;
 buffer[4244] = 16'h6023;
 buffer[4245] = 16'h6103;
 buffer[4246] = 16'h808C;
 buffer[4247] = 16'h6600;
 buffer[4248] = 16'h6023;
 buffer[4249] = 16'h6103;
 buffer[4250] = 16'h808D;
 buffer[4251] = 16'h6600;
 buffer[4252] = 16'h6023;
 buffer[4253] = 16'h6103;
 buffer[4254] = 16'h808E;
 buffer[4255] = 16'h6600;
 buffer[4256] = 16'h6023;
 buffer[4257] = 16'h6103;
 buffer[4258] = 16'h8001;
 buffer[4259] = 16'h808B;
 buffer[4260] = 16'h6600;
 buffer[4261] = 16'h6023;
 buffer[4262] = 16'h710F;
 buffer[4263] = 16'h211A;
 buffer[4264] = 16'h7404;
 buffer[4265] = 16'h7570;
 buffer[4266] = 16'h0021;
 buffer[4267] = 16'h80EA;
 buffer[4268] = 16'h6600;
 buffer[4269] = 16'h6C00;
 buffer[4270] = 16'h6010;
 buffer[4271] = 16'h30AB;
 buffer[4272] = 16'h80EA;
 buffer[4273] = 16'h6600;
 buffer[4274] = 16'h6023;
 buffer[4275] = 16'h710F;
 buffer[4276] = 16'h2150;
 buffer[4277] = 16'h7406;
 buffer[4278] = 16'h7570;
 buffer[4279] = 16'h7978;
 buffer[4280] = 16'h0021;
 buffer[4281] = 16'h80EE;
 buffer[4282] = 16'h6600;
 buffer[4283] = 16'h6023;
 buffer[4284] = 16'h6103;
 buffer[4285] = 16'h80EF;
 buffer[4286] = 16'h6600;
 buffer[4287] = 16'h6023;
 buffer[4288] = 16'h6103;
 buffer[4289] = 16'h8001;
 buffer[4290] = 16'h10AB;
 buffer[4291] = 16'h216A;
 buffer[4292] = 16'h740E;
 buffer[4293] = 16'h7570;
 buffer[4294] = 16'h6F66;
 buffer[4295] = 16'h6572;
 buffer[4296] = 16'h7267;
 buffer[4297] = 16'h756F;
 buffer[4298] = 16'h646E;
 buffer[4299] = 16'h0021;
 buffer[4300] = 16'h80EB;
 buffer[4301] = 16'h6600;
 buffer[4302] = 16'h6023;
 buffer[4303] = 16'h710F;
 buffer[4304] = 16'h2188;
 buffer[4305] = 16'h740E;
 buffer[4306] = 16'h7570;
 buffer[4307] = 16'h6162;
 buffer[4308] = 16'h6B63;
 buffer[4309] = 16'h7267;
 buffer[4310] = 16'h756F;
 buffer[4311] = 16'h646E;
 buffer[4312] = 16'h0021;
 buffer[4313] = 16'h80EC;
 buffer[4314] = 16'h6600;
 buffer[4315] = 16'h6023;
 buffer[4316] = 16'h710F;
 buffer[4317] = 16'h21A2;
 buffer[4318] = 16'h7407;
 buffer[4319] = 16'h7570;
 buffer[4320] = 16'h6D65;
 buffer[4321] = 16'h7469;
 buffer[4322] = 16'h80ED;
 buffer[4323] = 16'h6600;
 buffer[4324] = 16'h6023;
 buffer[4325] = 16'h6103;
 buffer[4326] = 16'h8002;
 buffer[4327] = 16'h10AB;
 buffer[4328] = 16'h21BC;
 buffer[4329] = 16'h7406;
 buffer[4330] = 16'h7570;
 buffer[4331] = 16'h7363;
 buffer[4332] = 16'h0021;
 buffer[4333] = 16'h8003;
 buffer[4334] = 16'h10AB;
 buffer[4335] = 16'h21D2;
 buffer[4336] = 16'h7408;
 buffer[4337] = 16'h7570;
 buffer[4338] = 16'h7073;
 buffer[4339] = 16'h6361;
 buffer[4340] = 16'h0065;
 buffer[4341] = 16'h4353;
 buffer[4342] = 16'h10E2;
 buffer[4343] = 16'h21E0;
 buffer[4344] = 16'h7409;
 buffer[4345] = 16'h7570;
 buffer[4346] = 16'h7073;
 buffer[4347] = 16'h6361;
 buffer[4348] = 16'h7365;
 buffer[4349] = 16'h8000;
 buffer[4350] = 16'h6E13;
 buffer[4351] = 16'h6147;
 buffer[4352] = 16'h1102;
 buffer[4353] = 16'h50F5;
 buffer[4354] = 16'h6B81;
 buffer[4355] = 16'h3108;
 buffer[4356] = 16'h6B8D;
 buffer[4357] = 16'h6A00;
 buffer[4358] = 16'h6147;
 buffer[4359] = 16'h1101;
 buffer[4360] = 16'h6B8D;
 buffer[4361] = 16'h710F;
 buffer[4362] = 16'h21F0;
 buffer[4363] = 16'h7407;
 buffer[4364] = 16'h7570;
 buffer[4365] = 16'h7974;
 buffer[4366] = 16'h6570;
 buffer[4367] = 16'h6147;
 buffer[4368] = 16'h1113;
 buffer[4369] = 16'h4383;
 buffer[4370] = 16'h50E2;
 buffer[4371] = 16'h6B81;
 buffer[4372] = 16'h3119;
 buffer[4373] = 16'h6B8D;
 buffer[4374] = 16'h6A00;
 buffer[4375] = 16'h6147;
 buffer[4376] = 16'h1111;
 buffer[4377] = 16'h6B8D;
 buffer[4378] = 16'h6103;
 buffer[4379] = 16'h710F;
 buffer[4380] = 16'h2216;
 buffer[4381] = 16'h7405;
 buffer[4382] = 16'h7570;
 buffer[4383] = 16'h242E;
 buffer[4384] = 16'h4383;
 buffer[4385] = 16'h110F;
 buffer[4386] = 16'h223A;
 buffer[4387] = 16'h7405;
 buffer[4388] = 16'h7570;
 buffer[4389] = 16'h722E;
 buffer[4390] = 16'h6147;
 buffer[4391] = 16'h441E;
 buffer[4392] = 16'h6B8D;
 buffer[4393] = 16'h6181;
 buffer[4394] = 16'h42A1;
 buffer[4395] = 16'h50FD;
 buffer[4396] = 16'h110F;
 buffer[4397] = 16'h2246;
 buffer[4398] = 16'h7406;
 buffer[4399] = 16'h7570;
 buffer[4400] = 16'h2E75;
 buffer[4401] = 16'h0072;
 buffer[4402] = 16'h6147;
 buffer[4403] = 16'h43EB;
 buffer[4404] = 16'h4404;
 buffer[4405] = 16'h4415;
 buffer[4406] = 16'h6B8D;
 buffer[4407] = 16'h6181;
 buffer[4408] = 16'h42A1;
 buffer[4409] = 16'h50FD;
 buffer[4410] = 16'h110F;
 buffer[4411] = 16'h225C;
 buffer[4412] = 16'h7405;
 buffer[4413] = 16'h7570;
 buffer[4414] = 16'h2E75;
 buffer[4415] = 16'h43EB;
 buffer[4416] = 16'h4404;
 buffer[4417] = 16'h4415;
 buffer[4418] = 16'h50F5;
 buffer[4419] = 16'h110F;
 buffer[4420] = 16'h2278;
 buffer[4421] = 16'h7404;
 buffer[4422] = 16'h7570;
 buffer[4423] = 16'h002E;
 buffer[4424] = 16'hFE80;
 buffer[4425] = 16'h6C00;
 buffer[4426] = 16'h800A;
 buffer[4427] = 16'h6503;
 buffer[4428] = 16'h314E;
 buffer[4429] = 16'h113F;
 buffer[4430] = 16'h441E;
 buffer[4431] = 16'h50F5;
 buffer[4432] = 16'h110F;
 buffer[4433] = 16'h228A;
 buffer[4434] = 16'h7405;
 buffer[4435] = 16'h7570;
 buffer[4436] = 16'h232E;
 buffer[4437] = 16'hFE80;
 buffer[4438] = 16'h6C00;
 buffer[4439] = 16'h6180;
 buffer[4440] = 16'h4432;
 buffer[4441] = 16'h5148;
 buffer[4442] = 16'hFE80;
 buffer[4443] = 16'h6023;
 buffer[4444] = 16'h710F;
 buffer[4445] = 16'h22A4;
 buffer[4446] = 16'h7406;
 buffer[4447] = 16'h7570;
 buffer[4448] = 16'h2E75;
 buffer[4449] = 16'h0023;
 buffer[4450] = 16'hFE80;
 buffer[4451] = 16'h6C00;
 buffer[4452] = 16'h6180;
 buffer[4453] = 16'h4432;
 buffer[4454] = 16'h43EB;
 buffer[4455] = 16'h4404;
 buffer[4456] = 16'h4415;
 buffer[4457] = 16'h50F5;
 buffer[4458] = 16'h510F;
 buffer[4459] = 16'hFE80;
 buffer[4460] = 16'h6023;
 buffer[4461] = 16'h710F;
 buffer[4462] = 16'h22BC;
 buffer[4463] = 16'h7407;
 buffer[4464] = 16'h7570;
 buffer[4465] = 16'h2E75;
 buffer[4466] = 16'h2372;
 buffer[4467] = 16'hFE80;
 buffer[4468] = 16'h6C00;
 buffer[4469] = 16'h427E;
 buffer[4470] = 16'h427E;
 buffer[4471] = 16'h4432;
 buffer[4472] = 16'h6147;
 buffer[4473] = 16'h43EB;
 buffer[4474] = 16'h4404;
 buffer[4475] = 16'h4415;
 buffer[4476] = 16'h6B8D;
 buffer[4477] = 16'h6181;
 buffer[4478] = 16'h42A1;
 buffer[4479] = 16'h50FD;
 buffer[4480] = 16'h510F;
 buffer[4481] = 16'hFE80;
 buffer[4482] = 16'h6023;
 buffer[4483] = 16'h710F;
 buffer[4484] = 16'h22DE;
 buffer[4485] = 16'h7406;
 buffer[4486] = 16'h7570;
 buffer[4487] = 16'h722E;
 buffer[4488] = 16'h0023;
 buffer[4489] = 16'hFE80;
 buffer[4490] = 16'h6C00;
 buffer[4491] = 16'h427E;
 buffer[4492] = 16'h427E;
 buffer[4493] = 16'h4432;
 buffer[4494] = 16'h6147;
 buffer[4495] = 16'h441E;
 buffer[4496] = 16'h6B8D;
 buffer[4497] = 16'h6181;
 buffer[4498] = 16'h42A1;
 buffer[4499] = 16'h50FD;
 buffer[4500] = 16'h510F;
 buffer[4501] = 16'hFE80;
 buffer[4502] = 16'h6023;
 buffer[4503] = 16'h710F;
 buffer[4504] = 16'h230A;
 buffer[4505] = 16'h7407;
 buffer[4506] = 16'h746D;
 buffer[4507] = 16'h6C69;
 buffer[4508] = 16'h2165;
 buffer[4509] = 16'h8069;
 buffer[4510] = 16'h6600;
 buffer[4511] = 16'h6023;
 buffer[4512] = 16'h6103;
 buffer[4513] = 16'h8010;
 buffer[4514] = 16'h6A00;
 buffer[4515] = 16'h6081;
 buffer[4516] = 16'h8068;
 buffer[4517] = 16'h6600;
 buffer[4518] = 16'h6023;
 buffer[4519] = 16'h6103;
 buffer[4520] = 16'h6180;
 buffer[4521] = 16'h8067;
 buffer[4522] = 16'h6600;
 buffer[4523] = 16'h6023;
 buffer[4524] = 16'h6103;
 buffer[4525] = 16'h6081;
 buffer[4526] = 16'h6010;
 buffer[4527] = 16'h31A2;
 buffer[4528] = 16'h710F;
 buffer[4529] = 16'h2332;
 buffer[4530] = 16'h7403;
 buffer[4531] = 16'h216D;
 buffer[4532] = 16'h806B;
 buffer[4533] = 16'h6600;
 buffer[4534] = 16'h6023;
 buffer[4535] = 16'h6103;
 buffer[4536] = 16'h806C;
 buffer[4537] = 16'h6600;
 buffer[4538] = 16'h6023;
 buffer[4539] = 16'h6103;
 buffer[4540] = 16'h806D;
 buffer[4541] = 16'h6600;
 buffer[4542] = 16'h6023;
 buffer[4543] = 16'h6103;
 buffer[4544] = 16'h806E;
 buffer[4545] = 16'h6600;
 buffer[4546] = 16'h6023;
 buffer[4547] = 16'h6103;
 buffer[4548] = 16'h806F;
 buffer[4549] = 16'h6600;
 buffer[4550] = 16'h6023;
 buffer[4551] = 16'h6103;
 buffer[4552] = 16'h8001;
 buffer[4553] = 16'h806A;
 buffer[4554] = 16'h6600;
 buffer[4555] = 16'h6023;
 buffer[4556] = 16'h710F;
 buffer[4557] = 16'h2364;
 buffer[4558] = 16'h7407;
 buffer[4559] = 16'h6D6D;
 buffer[4560] = 16'h766F;
 buffer[4561] = 16'h2165;
 buffer[4562] = 16'h8065;
 buffer[4563] = 16'h6600;
 buffer[4564] = 16'h6C00;
 buffer[4565] = 16'h6010;
 buffer[4566] = 16'h31D2;
 buffer[4567] = 16'h8066;
 buffer[4568] = 16'h6600;
 buffer[4569] = 16'h6023;
 buffer[4570] = 16'h710F;
 buffer[4571] = 16'h239C;
 buffer[4572] = 16'h7405;
 buffer[4573] = 16'h636D;
 buffer[4574] = 16'h2173;
 buffer[4575] = 16'h8065;
 buffer[4576] = 16'h6600;
 buffer[4577] = 16'h6C00;
 buffer[4578] = 16'h6010;
 buffer[4579] = 16'h31DF;
 buffer[4580] = 16'h8009;
 buffer[4581] = 16'h8066;
 buffer[4582] = 16'h6600;
 buffer[4583] = 16'h6023;
 buffer[4584] = 16'h710F;
 buffer[4585] = 16'h23B8;
 buffer[4586] = 16'h740D;
 buffer[4587] = 16'h7265;
 buffer[4588] = 16'h696D;
 buffer[4589] = 16'h616E;
 buffer[4590] = 16'h736C;
 buffer[4591] = 16'h6F68;
 buffer[4592] = 16'h2177;
 buffer[4593] = 16'h8001;
 buffer[4594] = 16'h80DE;
 buffer[4595] = 16'h6600;
 buffer[4596] = 16'h6023;
 buffer[4597] = 16'h710F;
 buffer[4598] = 16'h23D4;
 buffer[4599] = 16'h740D;
 buffer[4600] = 16'h7265;
 buffer[4601] = 16'h696D;
 buffer[4602] = 16'h616E;
 buffer[4603] = 16'h686C;
 buffer[4604] = 16'h6469;
 buffer[4605] = 16'h2165;
 buffer[4606] = 16'h8000;
 buffer[4607] = 16'h80DE;
 buffer[4608] = 16'h6600;
 buffer[4609] = 16'h6023;
 buffer[4610] = 16'h710F;
end

endmodule

module M_main (
in_btns,
in_uart_rx,
out_leds,
out_gpdi_dp,
out_gpdi_dn,
out_uart_tx,
out_audio_l,
out_audio_r,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [6:0] in_btns;
input  [0:0] in_uart_rx;
output  [7:0] out_leds;
output  [3:0] out_gpdi_dp;
output  [3:0] out_gpdi_dn;
output  [0:0] out_uart_tx;
output  [3:0] out_audio_l;
output  [3:0] out_audio_r;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = _w_clk_gen_clkout0;
wire _w_vga_rstcond_out;
wire _w_clk_gen_clkout0;
wire _w_clk_gen_clkout1;
wire _w_clk_gen_locked;
wire  [9:0] _w_video_x;
wire  [9:0] _w_video_y;
wire  [0:0] _w_video_active;
wire  [0:0] _w_video_vblank;
wire  [3:0] _w_video_gpdi_dp;
wire  [3:0] _w_video_gpdi_dn;
wire  [15:0] _w_ALU_newStackTop;
wire _w_ALU_done;
wire  [15:0] _w_CALLBRANCH_newStackTop;
wire  [12:0] _w_CALLBRANCH_newPC;
wire  [7:0] _w_CALLBRANCH_newDSP;
wire  [7:0] _w_CALLBRANCH_newRSP;
wire _w_CALLBRANCH_done;
wire  [7:0] _w_IO_Map_leds;
wire  [0:0] _w_IO_Map_uart_tx;
wire  [3:0] _w_IO_Map_audio_l;
wire  [3:0] _w_IO_Map_audio_r;
wire  [7:0] _w_IO_Map_video_r;
wire  [7:0] _w_IO_Map_video_g;
wire  [7:0] _w_IO_Map_video_b;
wire  [15:0] _w_IO_Map_readData;
wire _w_IO_Map_done;
wire  [15:0] _w_mem_dstack_rdata0;
wire  [15:0] _w_mem_rstack_rdata0;
wire  [15:0] _w_mem_ram_rdata0;
wire  [15:0] _w_immediate;
wire  [0:0] _w_is_alu;
wire  [0:0] _w_is_call;
wire  [0:0] _w_is_lit;
wire  [0:0] _w_is_n2memt;
wire  [1:0] _w_is_callbranchalu;
wire  [0:0] _w_dstackWrite;
wire  [0:0] _w_rstackWrite;
wire  [7:0] _w_ddelta;
wire  [7:0] _w_rdelta;
wire  [12:0] _w_pcPlusOne;
wire  [12:0] _w_callBranchAddress;
wire  [15:0] _w_stackNext;
wire  [15:0] _w_rStackTop;
wire  [15:0] _w_IOmemoryRead;
wire  [15:0] _w_RAMmemoryRead;

reg  [15:0] _d_instruction;
reg  [15:0] _q_instruction;
reg  [12:0] _d_pc;
reg  [12:0] _q_pc;
reg  [12:0] _d_newPC;
reg  [12:0] _q_newPC;
reg  [7:0] _d_dstack_addr0;
reg  [7:0] _q_dstack_addr0;
reg  [0:0] _d_dstack_wenable1;
reg  [0:0] _q_dstack_wenable1;
reg  [15:0] _d_dstack_wdata1;
reg  [15:0] _q_dstack_wdata1;
reg  [7:0] _d_dstack_addr1;
reg  [7:0] _q_dstack_addr1;
reg  [15:0] _d_stackTop;
reg  [15:0] _q_stackTop;
reg  [7:0] _d_dsp;
reg  [7:0] _q_dsp;
reg  [7:0] _d_newDSP;
reg  [7:0] _q_newDSP;
reg  [15:0] _d_newStackTop;
reg  [15:0] _q_newStackTop;
reg  [7:0] _d_rstack_addr0;
reg  [7:0] _q_rstack_addr0;
reg  [0:0] _d_rstack_wenable1;
reg  [0:0] _q_rstack_wenable1;
reg  [15:0] _d_rstack_wdata1;
reg  [15:0] _q_rstack_wdata1;
reg  [7:0] _d_rstack_addr1;
reg  [7:0] _q_rstack_addr1;
reg  [7:0] _d_rsp;
reg  [7:0] _q_rsp;
reg  [7:0] _d_newRSP;
reg  [7:0] _q_newRSP;
reg  [15:0] _d_rstackWData;
reg  [15:0] _q_rstackWData;
reg  [13:0] _d_ram_addr0;
reg  [13:0] _q_ram_addr0;
reg  [0:0] _d_ram_wenable1;
reg  [0:0] _q_ram_wenable1;
reg  [15:0] _d_ram_wdata1;
reg  [15:0] _q_ram_wdata1;
reg  [13:0] _d_ram_addr1;
reg  [13:0] _q_ram_addr1;
reg  [0:0] _d_IO_Map_memoryWrite,_q_IO_Map_memoryWrite;
reg  [0:0] _d_IO_Map_memoryRead,_q_IO_Map_memoryRead;
reg  [2:0] _d_index,_q_index;
reg  _ALU_run;
reg  _CALLBRANCH_run;
reg  _IO_Map_run;
assign out_leds = _w_IO_Map_leds;
assign out_gpdi_dp = _w_video_gpdi_dp;
assign out_gpdi_dn = _w_video_gpdi_dn;
assign out_uart_tx = _w_IO_Map_uart_tx;
assign out_audio_l = _w_IO_Map_audio_l;
assign out_audio_r = _w_IO_Map_audio_r;
assign out_done = (_q_index == 7);

always @(posedge _w_clk_gen_clkout0) begin
  if (reset || !in_run) begin
_q_pc <= 0;
_q_dstack_addr0 <= 0;
_q_dstack_wenable1 <= 0;
_q_dstack_wdata1 <= 0;
_q_dstack_addr1 <= 0;
_q_stackTop <= 0;
_q_dsp <= 0;
_q_rstack_addr0 <= 0;
_q_rstack_wenable1 <= 0;
_q_rstack_wdata1 <= 0;
_q_rstack_addr1 <= 0;
_q_rsp <= 0;
_q_ram_addr0 <= 0;
_q_ram_wenable1 <= 0;
_q_ram_wdata1 <= 0;
_q_ram_addr1 <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_instruction <= _d_instruction;
_q_pc <= _d_pc;
_q_newPC <= _d_newPC;
_q_dstack_addr0 <= _d_dstack_addr0;
_q_dstack_wenable1 <= _d_dstack_wenable1;
_q_dstack_wdata1 <= _d_dstack_wdata1;
_q_dstack_addr1 <= _d_dstack_addr1;
_q_stackTop <= _d_stackTop;
_q_dsp <= _d_dsp;
_q_newDSP <= _d_newDSP;
_q_newStackTop <= _d_newStackTop;
_q_rstack_addr0 <= _d_rstack_addr0;
_q_rstack_wenable1 <= _d_rstack_wenable1;
_q_rstack_wdata1 <= _d_rstack_wdata1;
_q_rstack_addr1 <= _d_rstack_addr1;
_q_rsp <= _d_rsp;
_q_newRSP <= _d_newRSP;
_q_rstackWData <= _d_rstackWData;
_q_ram_addr0 <= _d_ram_addr0;
_q_ram_wenable1 <= _d_ram_wenable1;
_q_ram_wdata1 <= _d_ram_wdata1;
_q_ram_addr1 <= _d_ram_addr1;
_q_index <= _d_index;
  end
_q_IO_Map_memoryWrite <= _d_IO_Map_memoryWrite;
_q_IO_Map_memoryRead <= _d_IO_Map_memoryRead;
end


reset_conditioner _vga_rstcond (
.rcclk(_w_clk_gen_clkout1),
.in(reset),
.out(_w_vga_rstcond_out)
);

ulx3s_clk_50_25 _clk_gen (
.clkin(clock),
.clkout0(_w_clk_gen_clkout0),
.clkout1(_w_clk_gen_clkout1),
.locked(_w_clk_gen_locked)
);
M_hdmi video (
.in_red(_w_IO_Map_video_r),
.in_green(_w_IO_Map_video_g),
.in_blue(_w_IO_Map_video_b),
.out_x(_w_video_x),
.out_y(_w_video_y),
.out_active(_w_video_active),
.out_vblank(_w_video_vblank),
.out_gpdi_dp(_w_video_gpdi_dp),
.out_gpdi_dn(_w_video_gpdi_dn),
.reset(reset),
.clock(clock)
);
M_j1eforthplusALU ALU (
.in_instruction(_d_instruction),
.in_dsp(_d_dsp),
.in_rsp(_d_rsp),
.in_stackTop(_d_stackTop),
.in_stackNext(_w_stackNext),
.in_rStackTop(_w_rStackTop),
.in_IOmemoryRead(_w_IOmemoryRead),
.in_RAMmemoryRead(_w_RAMmemoryRead),
.out_newStackTop(_w_ALU_newStackTop),
.out_done(_w_ALU_done),
.in_run(_ALU_run),
.reset(reset),
.clock(_w_clk_gen_clkout0)
);
M_j1eforthcallbranch CALLBRANCH (
.in_is_callbranchalu(_w_is_callbranchalu),
.in_stackTop(_d_stackTop),
.in_stackNext(_w_stackNext),
.in_callBranchAddress(_w_callBranchAddress),
.in_pcPlusOne(_w_pcPlusOne),
.in_dsp(_d_dsp),
.in_rsp(_d_rsp),
.out_newStackTop(_w_CALLBRANCH_newStackTop),
.out_newPC(_w_CALLBRANCH_newPC),
.out_newDSP(_w_CALLBRANCH_newDSP),
.out_newRSP(_w_CALLBRANCH_newRSP),
.out_done(_w_CALLBRANCH_done),
.in_run(_CALLBRANCH_run),
.reset(reset),
.clock(_w_clk_gen_clkout0)
);
M_memmap_io IO_Map (
.in_btns(in_btns),
.in_uart_rx(in_uart_rx),
.in_vblank(_w_video_vblank),
.in_pix_active(_w_video_active),
.in_pix_x(_w_video_x),
.in_pix_y(_w_video_y),
.in_clock_50mhz(_w_clk_gen_clkout0),
.in_clock_25mhz(clock),
.in_video_clock(_w_clk_gen_clkout1),
.in_video_reset(_w_vga_rstcond_out),
.in_memoryAddress(_d_stackTop),
.in_writeData(_w_stackNext),
.in_memoryWrite(_d_IO_Map_memoryWrite),
.in_memoryRead(_d_IO_Map_memoryRead),
.out_leds(_w_IO_Map_leds),
.out_uart_tx(_w_IO_Map_uart_tx),
.out_audio_l(_w_IO_Map_audio_l),
.out_audio_r(_w_IO_Map_audio_r),
.out_video_r(_w_IO_Map_video_r),
.out_video_g(_w_IO_Map_video_g),
.out_video_b(_w_IO_Map_video_b),
.out_readData(_w_IO_Map_readData),
.out_done(_w_IO_Map_done),
.in_run(_IO_Map_run),
.reset(reset),
.clock(_w_clk_gen_clkout0)
);

M_main_mem_dstack __mem__dstack(
.clock0(_w_clk_gen_clkout0),
.clock1(_w_clk_gen_clkout0),
.in_dstack_addr0(_d_dstack_addr0),
.in_dstack_wenable1(_d_dstack_wenable1),
.in_dstack_wdata1(_d_dstack_wdata1),
.in_dstack_addr1(_d_dstack_addr1),
.out_dstack_rdata0(_w_mem_dstack_rdata0)
);
M_main_mem_rstack __mem__rstack(
.clock0(_w_clk_gen_clkout0),
.clock1(_w_clk_gen_clkout0),
.in_rstack_addr0(_d_rstack_addr0),
.in_rstack_wenable1(_d_rstack_wenable1),
.in_rstack_wdata1(_d_rstack_wdata1),
.in_rstack_addr1(_d_rstack_addr1),
.out_rstack_rdata0(_w_mem_rstack_rdata0)
);
M_main_mem_ram __mem__ram(
.clock0(_w_clk_gen_clkout0),
.clock1(_w_clk_gen_clkout0),
.in_ram_addr0(_d_ram_addr0),
.in_ram_wenable1(_d_ram_wenable1),
.in_ram_wdata1(_d_ram_wdata1),
.in_ram_addr1(_d_ram_addr1),
.out_ram_rdata0(_w_mem_ram_rdata0)
);

assign _w_rStackTop = _w_mem_rstack_rdata0;
assign _w_immediate = (_d_instruction[0+:15]);
assign _w_is_alu = (_d_instruction[13+:3]==3'b011);
assign _w_is_lit = _d_instruction[15+:1];
assign _w_is_call = (_d_instruction[13+:3]==3'b010);
assign _w_RAMmemoryRead = _w_mem_ram_rdata0;
assign _w_IOmemoryRead = _w_IO_Map_readData;
assign _w_ddelta = {{7{_d_instruction[1+:1]}},_d_instruction[0+:1]};
assign _w_callBranchAddress = _d_instruction[0+:13];
assign _w_is_n2memt = _w_is_alu&&_d_instruction[5+:1];
assign _w_is_callbranchalu = _d_instruction[13+:2];
assign _w_dstackWrite = (_w_is_lit|(_w_is_alu&_d_instruction[7+:1]));
assign _w_rdelta = {{7{_d_instruction[3+:1]}},_d_instruction[2+:1]};
assign _w_pcPlusOne = _d_pc+1;
assign _w_rstackWrite = (_w_is_call|(_w_is_alu&_d_instruction[6+:1]));
assign _w_stackNext = _w_mem_dstack_rdata0;

always @* begin
_d_instruction = _q_instruction;
_d_pc = _q_pc;
_d_newPC = _q_newPC;
_d_dstack_addr0 = _q_dstack_addr0;
_d_dstack_wenable1 = _q_dstack_wenable1;
_d_dstack_wdata1 = _q_dstack_wdata1;
_d_dstack_addr1 = _q_dstack_addr1;
_d_stackTop = _q_stackTop;
_d_dsp = _q_dsp;
_d_newDSP = _q_newDSP;
_d_newStackTop = _q_newStackTop;
_d_rstack_addr0 = _q_rstack_addr0;
_d_rstack_wenable1 = _q_rstack_wenable1;
_d_rstack_wdata1 = _q_rstack_wdata1;
_d_rstack_addr1 = _q_rstack_addr1;
_d_rsp = _q_rsp;
_d_newRSP = _q_newRSP;
_d_rstackWData = _q_rstackWData;
_d_ram_addr0 = _q_ram_addr0;
_d_ram_wenable1 = _q_ram_wenable1;
_d_ram_wdata1 = _q_ram_wdata1;
_d_ram_addr1 = _q_ram_addr1;
_d_IO_Map_memoryWrite = _q_IO_Map_memoryWrite;
_d_IO_Map_memoryRead = _q_IO_Map_memoryRead;
_d_index = _q_index;
_ALU_run = 1;
_CALLBRANCH_run = 1;
_IO_Map_run = 1;
// _always_pre
_d_ram_wenable1 = 1;
_d_dstack_addr0 = _q_dsp;
_d_dstack_wenable1 = 1;
_d_rstack_addr0 = _q_rsp;
_d_rstack_wenable1 = 1;
_d_IO_Map_memoryWrite = 0;
_d_IO_Map_memoryRead = 0;
_d_index = 7;
(* full_case *)
case (_q_index)
0: begin
// _top
// var inits
_d_pc = 0;
_d_dstack_addr0 = 0;
_d_dstack_wenable1 = 0;
_d_dstack_wdata1 = 0;
_d_dstack_addr1 = 0;
_d_stackTop = 0;
_d_dsp = 0;
_d_rstack_addr0 = 0;
_d_rstack_wenable1 = 0;
_d_rstack_wdata1 = 0;
_d_rstack_addr1 = 0;
_d_rsp = 0;
_d_ram_addr0 = 0;
_d_ram_wenable1 = 0;
_d_ram_wdata1 = 0;
_d_ram_addr1 = 0;
// --
_d_ram_addr1 = 16383;
_d_ram_wdata1 = 0;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
_d_ram_addr0 = _q_pc;
_d_index = 3;
end else begin
_d_index = 2;
end
end
3: begin
// __block_5
_d_instruction = _w_mem_ram_rdata0;
_d_ram_addr0 = _q_stackTop>>1;
_d_index = 4;
end
2: begin
// __block_3
_d_index = 7;
end
4: begin
// __block_6
if (_w_is_lit) begin
// __block_7
// __block_9
_d_newStackTop = _w_immediate;
_d_newPC = _w_pcPlusOne;
_d_newDSP = _q_dsp+1;
_d_newRSP = _q_rsp;
// __block_10
end else begin
// __block_8
// __block_11
  case (_q_instruction[13+:2])
  2'b11: begin
// __block_13_case
// __block_14
if (~_q_instruction[4+:1]&&(_q_instruction[8+:4]==4'b1100)&&_q_stackTop[15+:1]) begin
// __block_15
// __block_17
_d_IO_Map_memoryRead = 1;
// __block_18
end else begin
// __block_16
end
// __block_19
_d_newStackTop = _w_ALU_newStackTop;
_d_newDSP = _q_dsp+_w_ddelta;
_d_newRSP = _q_rsp+_w_rdelta;
_d_rstackWData = _q_stackTop;
_d_newPC = (_q_instruction[12+:1])?_w_rStackTop>>1:_w_pcPlusOne;
if (_w_is_n2memt&&~_q_stackTop[15+:1]) begin
// __block_20
// __block_22
_d_ram_addr1 = _q_stackTop>>1;
_d_ram_wdata1 = _w_stackNext;
// __block_23
end else begin
// __block_21
end
// __block_24
_d_IO_Map_memoryWrite = _w_is_n2memt&&(_q_stackTop[15+:1]);
// __block_25
  end
  default: begin
// __block_26_case
// __block_27
_d_newStackTop = _w_CALLBRANCH_newStackTop;
_d_newPC = _w_CALLBRANCH_newPC;
_d_newDSP = _w_CALLBRANCH_newDSP;
_d_newRSP = _w_CALLBRANCH_newRSP;
_d_rstackWData = _w_pcPlusOne<<1;
// __block_28
  end
endcase
// __block_12
// __block_29
end
// __block_30
_d_index = 5;
end
5: begin
// __block_31
if (_w_dstackWrite) begin
// __block_32
// __block_34
_d_dstack_addr1 = _q_newDSP;
_d_dstack_wdata1 = _q_stackTop;
// __block_35
end else begin
// __block_33
end
// __block_36
if (_w_rstackWrite) begin
// __block_37
// __block_39
_d_rstack_addr1 = _q_newRSP;
_d_rstack_wdata1 = _q_rstackWData;
// __block_40
end else begin
// __block_38
end
// __block_41
_d_dsp = _q_newDSP;
_d_pc = _q_newPC;
_d_stackTop = _q_newStackTop;
_d_rsp = _q_newRSP;
_d_index = 6;
end
6: begin
// __block_42
// __block_43
_d_index = 1;
end
7: begin // end of main
end
default: begin 
_d_index = 7;
 end
endcase
end
endmodule


module M_j1eforthplusALU (
in_instruction,
in_dsp,
in_rsp,
in_stackTop,
in_stackNext,
in_rStackTop,
in_IOmemoryRead,
in_RAMmemoryRead,
out_newStackTop,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [15:0] in_instruction;
input  [7:0] in_dsp;
input  [7:0] in_rsp;
input  [15:0] in_stackTop;
input  [15:0] in_stackNext;
input  [15:0] in_rStackTop;
input  [15:0] in_IOmemoryRead;
input  [15:0] in_RAMmemoryRead;
output  [15:0] out_newStackTop;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [15:0] _d_newStackTop,_q_newStackTop;
reg  [1:0] _d_index,_q_index;
assign out_newStackTop = _d_newStackTop;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_newStackTop <= _d_newStackTop;
_q_index <= _d_index;
  end
end




always @* begin
_d_newStackTop = _q_newStackTop;
_d_index = _q_index;
// _always_pre
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (in_instruction[4+:1])
  1'b0: begin
// __block_6_case
// __block_7
  case (in_instruction[8+:4])
  4'b0000: begin
// __block_9_case
// __block_10
_d_newStackTop = in_stackTop;
// __block_11
  end
  4'b0001: begin
// __block_12_case
// __block_13
_d_newStackTop = in_stackNext;
// __block_14
  end
  4'b0010: begin
// __block_15_case
// __block_16
_d_newStackTop = in_stackTop+in_stackNext;
// __block_17
  end
  4'b0011: begin
// __block_18_case
// __block_19
_d_newStackTop = in_stackTop&in_stackNext;
// __block_20
  end
  4'b0100: begin
// __block_21_case
// __block_22
_d_newStackTop = in_stackTop|in_stackNext;
// __block_23
  end
  4'b0101: begin
// __block_24_case
// __block_25
_d_newStackTop = in_stackTop^in_stackNext;
// __block_26
  end
  4'b0110: begin
// __block_27_case
// __block_28
_d_newStackTop = ~in_stackTop;
// __block_29
  end
  4'b0111: begin
// __block_30_case
// __block_31
_d_newStackTop = {16{(in_stackNext==in_stackTop)}};
// __block_32
  end
  4'b1000: begin
// __block_33_case
// __block_34
_d_newStackTop = {16{($signed(in_stackNext)<$signed(in_stackTop))}};
// __block_35
  end
  4'b1001: begin
// __block_36_case
// __block_37
_d_newStackTop = in_stackNext>>in_stackTop[0+:4];
// __block_38
  end
  4'b1010: begin
// __block_39_case
// __block_40
_d_newStackTop = in_stackTop-1;
// __block_41
  end
  4'b1011: begin
// __block_42_case
// __block_43
_d_newStackTop = in_rStackTop;
// __block_44
  end
  4'b1100: begin
// __block_45_case
// __block_46
_d_newStackTop = in_stackTop[15+:1]?in_IOmemoryRead:in_RAMmemoryRead;
// __block_47
  end
  4'b1101: begin
// __block_48_case
// __block_49
_d_newStackTop = in_stackNext<<in_stackTop[0+:4];
// __block_50
  end
  4'b1110: begin
// __block_51_case
// __block_52
_d_newStackTop = {in_rsp,in_dsp};
// __block_53
  end
  4'b1111: begin
// __block_54_case
// __block_55
_d_newStackTop = {16{($unsigned(in_stackNext)<$unsigned(in_stackTop))}};
// __block_56
  end
endcase
// __block_8
// __block_57
  end
  1'b1: begin
// __block_58_case
// __block_59
  case (in_instruction[8+:4])
  4'b0000: begin
// __block_61_case
// __block_62
_d_newStackTop = {16{(in_stackTop==0)}};
// __block_63
  end
  4'b0001: begin
// __block_64_case
// __block_65
_d_newStackTop = {16{(in_stackTop!=0)}};
// __block_66
  end
  4'b0010: begin
// __block_67_case
// __block_68
_d_newStackTop = {16{(in_stackNext!=in_stackTop)}};
// __block_69
  end
  4'b0011: begin
// __block_70_case
// __block_71
_d_newStackTop = in_stackTop+1;
// __block_72
  end
  4'b0100: begin
// __block_73_case
// __block_74
_d_newStackTop = in_stackNext*in_stackTop;
// __block_75
  end
  4'b0101: begin
// __block_76_case
// __block_77
_d_newStackTop = in_stackTop<<1;
// __block_78
  end
  4'b0110: begin
// __block_79_case
// __block_80
_d_newStackTop = -in_stackTop;
// __block_81
  end
  4'b0111: begin
// __block_82_case
// __block_83
_d_newStackTop = {in_stackTop[15+:1],in_stackTop[1+:15]};
// __block_84
  end
  4'b1000: begin
// __block_85_case
// __block_86
_d_newStackTop = in_stackNext-in_stackTop;
// __block_87
  end
  4'b1001: begin
// __block_88_case
// __block_89
_d_newStackTop = {16{($signed(in_stackTop)<$signed(0))}};
// __block_90
  end
  4'b1010: begin
// __block_91_case
// __block_92
_d_newStackTop = {16{($signed(in_stackTop)>$signed(0))}};
// __block_93
  end
  4'b1011: begin
// __block_94_case
// __block_95
_d_newStackTop = {16{($signed(in_stackNext)>$signed(in_stackTop))}};
// __block_96
  end
  4'b1100: begin
// __block_97_case
// __block_98
_d_newStackTop = {16{($signed(in_stackNext)>=$signed(in_stackTop))}};
// __block_99
  end
  4'b1101: begin
// __block_100_case
// __block_101
_d_newStackTop = ($signed(in_stackTop)<$signed(0))?-in_stackTop:in_stackTop;
// __block_102
  end
  4'b1110: begin
// __block_103_case
// __block_104
_d_newStackTop = ($signed(in_stackNext)>$signed(in_stackTop))?in_stackNext:in_stackTop;
// __block_105
  end
  4'b1111: begin
// __block_106_case
// __block_107
_d_newStackTop = ($signed(in_stackNext)<$signed(in_stackTop))?in_stackNext:in_stackTop;
// __block_108
  end
endcase
// __block_60
// __block_109
  end
endcase
// __block_5
// __block_110
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of j1eforthplusALU
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_j1eforthcallbranch (
in_is_callbranchalu,
in_stackTop,
in_stackNext,
in_callBranchAddress,
in_pcPlusOne,
in_dsp,
in_rsp,
out_newStackTop,
out_newPC,
out_newDSP,
out_newRSP,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [1:0] in_is_callbranchalu;
input  [15:0] in_stackTop;
input  [15:0] in_stackNext;
input  [12:0] in_callBranchAddress;
input  [12:0] in_pcPlusOne;
input  [7:0] in_dsp;
input  [7:0] in_rsp;
output  [15:0] out_newStackTop;
output  [12:0] out_newPC;
output  [7:0] out_newDSP;
output  [7:0] out_newRSP;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg  [15:0] _d_newStackTop,_q_newStackTop;
reg  [12:0] _d_newPC,_q_newPC;
reg  [7:0] _d_newDSP,_q_newDSP;
reg  [7:0] _d_newRSP,_q_newRSP;
reg  [1:0] _d_index,_q_index;
assign out_newStackTop = _d_newStackTop;
assign out_newPC = _d_newPC;
assign out_newDSP = _d_newDSP;
assign out_newRSP = _d_newRSP;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_newStackTop <= _d_newStackTop;
_q_newPC <= _d_newPC;
_q_newDSP <= _d_newDSP;
_q_newRSP <= _d_newRSP;
_q_index <= _d_index;
  end
end




always @* begin
_d_newStackTop = _q_newStackTop;
_d_newPC = _q_newPC;
_d_newDSP = _q_newDSP;
_d_newRSP = _q_newRSP;
_d_index = _q_index;
// _always_pre
_d_index = 3;
(* full_case *)
case (_q_index)
0: begin
// _top
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (in_is_callbranchalu)
  2'b00: begin
// __block_6_case
// __block_7
_d_newStackTop = in_stackTop;
_d_newPC = in_callBranchAddress;
_d_newDSP = in_dsp;
_d_newRSP = in_rsp;
// __block_8
  end
  2'b01: begin
// __block_9_case
// __block_10
_d_newStackTop = in_stackNext;
_d_newPC = (in_stackTop==0)?in_callBranchAddress:in_pcPlusOne;
_d_newDSP = in_dsp-1;
_d_newRSP = in_rsp;
// __block_11
  end
  2'b10: begin
// __block_12_case
// __block_13
_d_newStackTop = in_stackTop;
_d_newPC = in_callBranchAddress;
_d_newDSP = in_dsp;
_d_newRSP = in_rsp+1;
// __block_14
  end
endcase
// __block_5
// __block_15
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of j1eforthcallbranch
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule

