`define DE10NANO 1

module Basic(
    // 50MHz clock input
    input clk,
    
    // uart via GPIO pins
    output tx,
    input rx,
    
    // Outputs to the 8 onboard LEDs
    output reg LED0,
    output reg LED1,
    output reg LED2,
    output reg LED3,
    output reg LED4,
    output reg LED5,
    output reg LED6,
    output reg LED7
    );

wire [7:0] __main_out_led;

reg [31:0] RST_d;
reg [31:0] RST_q;

reg ready = 0;

always @* begin
  RST_d = RST_q >> 1;
end

always @(posedge clk) begin
  if (ready) begin
    RST_q <= RST_d;
  end else begin
    ready <= 1;
    RST_q <= 32'b111111111111111111111111111111;
  end
end

wire reset_main;
assign reset_main = RST_q[0];
wire run_main;
assign run_main = 1'b1;


// Create 1hz (1 second counter)
reg [31:0] counter50mhz;
reg [15:0] counter1hz;
always @(posedge clk) begin
    if( counter50mhz == 50000000 ) begin
        counter1hz <= counter1hz + 1;
        counter50mhz <= 0;
    end else begin
        counter50mhz <= counter50mhz + 1;
    end
end 

// UART tx and rx
wire [7:0] uart_tx_data;
wire uart_tx_valid;
wire uart_tx_busy;
wire uart_tx_done;
wire [7:0] uart_rx_data;
wire uart_rx_valid;
wire uart_rx_ready;
wire uart_serial_tx;

//uart uart0(
//.clk(clk), // The master clock for this module
//.rst(reset_main), // Synchronous reset
//.rx(rx), // Incoming serial line
//.tx(tx), // Outgoing serial line
//.transmit(uart_tx_valid), // Signal to transmit
//.tx_byte(uart_tx_data), // Byte to transmit
//.received(uart_rx_valid), // Indicated that a byte has been received
//.rx_byte(uart_rx_data), // Byte received
//.is_receiving(), // Low when receive line is idle
//.is_transmitting(uart_tx_busy),// Low when transmit line is idle
//.recv_error() // Indicates error in receiving packet.
//);

// Want to interface to 115200 baud UART
// 50000000 / 115200 = 434 Clocks Per Bit.
parameter c_CLOCK_PERIOD_NS = 2;
parameter c_CLKS_PER_BIT    = 434;
parameter c_BIT_PERIOD      = 8600;

uart_rx #(.CLKS_PER_BIT(c_CLKS_PER_BIT)) UART_RX_INST
(.i_Clock(clk),
    .i_Rx_Serial(rx),
    .o_Rx_DV(uart_rx_valid),
    .o_Rx_Byte(uart_rx_data)
    );

uart_tx #(.CLKS_PER_BIT(c_CLKS_PER_BIT)) UART_TX_INST
(.i_Clock(clk),
    .i_Tx_DV(uart_tx_valid),
    .i_Tx_Byte(uart_tx_data),
    .o_Tx_Active(uart_tx_busy),
    .o_Tx_Serial(tx),
    .o_Tx_Done(uart_tx_done)
    );

M_main __main(
  .clock(clk),
  .reset(reset_main),
  .in_run(run_main),
  .out_led(__main_out_led),

  // UART
  .out_uart_tx_data( uart_tx_data ),
  .out_uart_tx_valid( uart_tx_valid ),
  .in_uart_tx_busy( uart_tx_busy ),

  .in_uart_rx_data( uart_rx_data ),
  .in_uart_rx_valid( uart_rx_valid ),
    
  .in_timer1hz ( counter1hz )
);

always @* begin
  LED0 = __main_out_led[0+:1];
  LED1 = __main_out_led[1+:1];
  LED2 = __main_out_led[2+:1];
  LED3 = __main_out_led[3+:1];
  LED4 = __main_out_led[4+:1];
  LED5 = __main_out_led[5+:1];
  LED6 = __main_out_led[6+:1];
  LED7 = __main_out_led[7+:1];
end

endmodule

module M_main_mem_dstack(
input                  [0:0] in_dstack_wenable,
input       [15:0]    in_dstack_wdata,
input                  [7:0]    in_dstack_addr,
output reg  [15:0]    out_dstack_rdata,
input                                      clock
);
reg  [15:0] buffer[255:0];
always @(posedge clock) begin
  if (in_dstack_wenable) begin
    buffer[in_dstack_addr] <= in_dstack_wdata;
  end
  out_dstack_rdata <= buffer[in_dstack_addr];
end

endmodule

module M_main_mem_rstack(
input                  [0:0] in_rstack_wenable,
input       [15:0]    in_rstack_wdata,
input                  [7:0]    in_rstack_addr,
output reg  [15:0]    out_rstack_rdata,
input                                      clock
);
reg  [15:0] buffer[255:0];
always @(posedge clock) begin
  if (in_rstack_wenable) begin
    buffer[in_rstack_addr] <= in_rstack_wdata;
  end
  out_rstack_rdata <= buffer[in_rstack_addr];
end

endmodule

module M_main_mem_rom(
input                  [11:0] in_rom_addr,
output reg  [15:0] out_rom_rdata,
input                                   clock
);
reg  [15:0] buffer[3609:0];
always @(posedge clock) begin
   out_rom_rdata <= buffer[in_rom_addr];
end
initial begin
 buffer[0] = 16'h0E02;
 buffer[1] = 16'h0010;
 buffer[2] = 16'h0000;
 buffer[3] = 16'h0000;
 buffer[4] = 16'h0000;
 buffer[5] = 16'h7F00;
 buffer[6] = 16'h1058;
 buffer[7] = 16'h1136;
 buffer[8] = 16'h0000;
 buffer[9] = 16'h0000;
 buffer[10] = 16'h0000;
 buffer[11] = 16'h0000;
 buffer[12] = 16'h0000;
 buffer[13] = 16'h0000;
 buffer[14] = 16'h0000;
 buffer[15] = 16'h0000;
 buffer[16] = 16'h0000;
 buffer[17] = 16'h0000;
 buffer[18] = 16'h0000;
 buffer[19] = 16'h0000;
 buffer[20] = 16'h0000;
 buffer[21] = 16'h0000;
 buffer[22] = 16'h0000;
 buffer[23] = 16'h1C34;
 buffer[24] = 16'h1BFE;
 buffer[25] = 16'h0952;
 buffer[26] = 16'h0964;
 buffer[27] = 16'h1BCA;
 buffer[28] = 16'h0E14;
 buffer[29] = 16'h0F00;
 buffer[30] = 16'h160C;
 buffer[31] = 16'h168E;
 buffer[32] = 16'h16B6;
 buffer[33] = 16'h1722;
 buffer[34] = 16'h0000;
 buffer[35] = 16'h0000;
 buffer[36] = 16'h0000;
 buffer[37] = 16'h0000;
 buffer[38] = 16'h0000;
 buffer[39] = 16'h0000;
 buffer[40] = 16'h0000;
 buffer[41] = 16'h0000;
 buffer[42] = 16'h0000;
 buffer[43] = 16'h0000;
 buffer[44] = 16'h0000;
 buffer[45] = 16'h0000;
 buffer[46] = 16'h0000;
 buffer[47] = 16'h0000;
 buffer[48] = 16'h0000;
 buffer[49] = 16'h0000;
 buffer[50] = 16'h0000;
 buffer[51] = 16'h0000;
 buffer[52] = 16'h0000;
 buffer[53] = 16'h0000;
 buffer[54] = 16'h0000;
 buffer[55] = 16'h0000;
 buffer[56] = 16'h0000;
 buffer[57] = 16'h0000;
 buffer[58] = 16'h0000;
 buffer[59] = 16'h0000;
 buffer[60] = 16'h0000;
 buffer[61] = 16'h0000;
 buffer[62] = 16'h0000;
 buffer[63] = 16'h0000;
 buffer[64] = 16'h6003;
 buffer[65] = 16'h6003;
 buffer[66] = 16'h6003;
 buffer[67] = 16'h6003;
 buffer[68] = 16'h6003;
 buffer[69] = 16'h6003;
 buffer[70] = 16'h6003;
 buffer[71] = 16'h6003;
 buffer[72] = 16'h6003;
 buffer[73] = 16'h6003;
 buffer[74] = 16'h6003;
 buffer[75] = 16'h6003;
 buffer[76] = 16'h6003;
 buffer[77] = 16'h6003;
 buffer[78] = 16'h6003;
 buffer[79] = 16'h710C;
 buffer[80] = 16'h6001;
 buffer[81] = 16'h6001;
 buffer[82] = 16'h6001;
 buffer[83] = 16'h6001;
 buffer[84] = 16'h6001;
 buffer[85] = 16'h6001;
 buffer[86] = 16'h6001;
 buffer[87] = 16'h6001;
 buffer[88] = 16'h6001;
 buffer[89] = 16'h6001;
 buffer[90] = 16'h6001;
 buffer[91] = 16'h6001;
 buffer[92] = 16'h6001;
 buffer[93] = 16'h6001;
 buffer[94] = 16'h6001;
 buffer[95] = 16'h700C;
 buffer[96] = 16'h6100;
 buffer[97] = 16'h700C;
 buffer[98] = 16'h404E;
 buffer[99] = 16'h005E;
 buffer[100] = 16'h404D;
 buffer[101] = 16'h005D;
 buffer[102] = 16'h404C;
 buffer[103] = 16'h005C;
 buffer[104] = 16'h404B;
 buffer[105] = 16'h005B;
 buffer[106] = 16'h404A;
 buffer[107] = 16'h005A;
 buffer[108] = 16'h4049;
 buffer[109] = 16'h0059;
 buffer[110] = 16'h4048;
 buffer[111] = 16'h0058;
 buffer[112] = 16'h4047;
 buffer[113] = 16'h0057;
 buffer[114] = 16'h4046;
 buffer[115] = 16'h0056;
 buffer[116] = 16'h4045;
 buffer[117] = 16'h0055;
 buffer[118] = 16'h4044;
 buffer[119] = 16'h0054;
 buffer[120] = 16'h4043;
 buffer[121] = 16'h0053;
 buffer[122] = 16'h4042;
 buffer[123] = 16'h0052;
 buffer[124] = 16'h4041;
 buffer[125] = 16'h0051;
 buffer[126] = 16'h4040;
 buffer[127] = 16'h0050;
 buffer[128] = 16'h700C;
 buffer[129] = 16'h0000;
 buffer[130] = 16'h0000;
 buffer[131] = 16'h0000;
 buffer[132] = 16'h0000;
 buffer[133] = 16'h0000;
 buffer[134] = 16'h0000;
 buffer[135] = 16'h0000;
 buffer[136] = 16'h0000;
 buffer[137] = 16'h0000;
 buffer[138] = 16'h0000;
 buffer[139] = 16'h0000;
 buffer[140] = 16'h0000;
 buffer[141] = 16'h0000;
 buffer[142] = 16'h0000;
 buffer[143] = 16'h0000;
 buffer[144] = 16'h0000;
 buffer[145] = 16'h0000;
 buffer[146] = 16'h0000;
 buffer[147] = 16'h0000;
 buffer[148] = 16'h0000;
 buffer[149] = 16'h0000;
 buffer[150] = 16'h0000;
 buffer[151] = 16'h0000;
 buffer[152] = 16'h0000;
 buffer[153] = 16'h0000;
 buffer[154] = 16'h0000;
 buffer[155] = 16'h0000;
 buffer[156] = 16'h0000;
 buffer[157] = 16'h0000;
 buffer[158] = 16'h0000;
 buffer[159] = 16'h0000;
 buffer[160] = 16'h0000;
 buffer[161] = 16'h0000;
 buffer[162] = 16'h0000;
 buffer[163] = 16'h0000;
 buffer[164] = 16'h0000;
 buffer[165] = 16'h0000;
 buffer[166] = 16'h0000;
 buffer[167] = 16'h0000;
 buffer[168] = 16'h0000;
 buffer[169] = 16'h0000;
 buffer[170] = 16'h0000;
 buffer[171] = 16'h0000;
 buffer[172] = 16'h0000;
 buffer[173] = 16'h0000;
 buffer[174] = 16'h0000;
 buffer[175] = 16'h0000;
 buffer[176] = 16'h0000;
 buffer[177] = 16'h0000;
 buffer[178] = 16'h0000;
 buffer[179] = 16'h0000;
 buffer[180] = 16'h0000;
 buffer[181] = 16'h0000;
 buffer[182] = 16'h0000;
 buffer[183] = 16'h0000;
 buffer[184] = 16'h0000;
 buffer[185] = 16'h0000;
 buffer[186] = 16'h0000;
 buffer[187] = 16'h0000;
 buffer[188] = 16'h0000;
 buffer[189] = 16'h0000;
 buffer[190] = 16'h0000;
 buffer[191] = 16'h0000;
 buffer[192] = 16'h0000;
 buffer[193] = 16'h6E04;
 buffer[194] = 16'h6F6F;
 buffer[195] = 16'h0070;
 buffer[196] = 16'h700C;
 buffer[197] = 16'h0182;
 buffer[198] = 16'h2B01;
 buffer[199] = 16'h720F;
 buffer[200] = 16'h018C;
 buffer[201] = 16'h7803;
 buffer[202] = 16'h726F;
 buffer[203] = 16'h750F;
 buffer[204] = 16'h0192;
 buffer[205] = 16'h6103;
 buffer[206] = 16'h646E;
 buffer[207] = 16'h730F;
 buffer[208] = 16'h019A;
 buffer[209] = 16'h6F02;
 buffer[210] = 16'h0072;
 buffer[211] = 16'h740F;
 buffer[212] = 16'h01A2;
 buffer[213] = 16'h6906;
 buffer[214] = 16'h766E;
 buffer[215] = 16'h7265;
 buffer[216] = 16'h0074;
 buffer[217] = 16'h760C;
 buffer[218] = 16'h01AA;
 buffer[219] = 16'h3D01;
 buffer[220] = 16'h770F;
 buffer[221] = 16'h01B6;
 buffer[222] = 16'h3C01;
 buffer[223] = 16'h780F;
 buffer[224] = 16'h01BC;
 buffer[225] = 16'h7502;
 buffer[226] = 16'h003C;
 buffer[227] = 16'h7F0F;
 buffer[228] = 16'h01C2;
 buffer[229] = 16'h7304;
 buffer[230] = 16'h6177;
 buffer[231] = 16'h0070;
 buffer[232] = 16'h718C;
 buffer[233] = 16'h01CA;
 buffer[234] = 16'h7502;
 buffer[235] = 16'h003E;
 buffer[236] = 16'h771F;
 buffer[237] = 16'h01D4;
 buffer[238] = 16'h6403;
 buffer[239] = 16'h7075;
 buffer[240] = 16'h708D;
 buffer[241] = 16'h01DC;
 buffer[242] = 16'h6404;
 buffer[243] = 16'h6F72;
 buffer[244] = 16'h0070;
 buffer[245] = 16'h710F;
 buffer[246] = 16'h01E4;
 buffer[247] = 16'h6F04;
 buffer[248] = 16'h6576;
 buffer[249] = 16'h0072;
 buffer[250] = 16'h718D;
 buffer[251] = 16'h01EE;
 buffer[252] = 16'h6E03;
 buffer[253] = 16'h7069;
 buffer[254] = 16'h700F;
 buffer[255] = 16'h01F8;
 buffer[256] = 16'h6C06;
 buffer[257] = 16'h6873;
 buffer[258] = 16'h6669;
 buffer[259] = 16'h0074;
 buffer[260] = 16'h7D0F;
 buffer[261] = 16'h0200;
 buffer[262] = 16'h7206;
 buffer[263] = 16'h6873;
 buffer[264] = 16'h6669;
 buffer[265] = 16'h0074;
 buffer[266] = 16'h790F;
 buffer[267] = 16'h020C;
 buffer[268] = 16'h3102;
 buffer[269] = 16'h002D;
 buffer[270] = 16'h7A0C;
 buffer[271] = 16'h0218;
 buffer[272] = 16'h3E42;
 buffer[273] = 16'h0072;
 buffer[274] = 16'h6B8D;
 buffer[275] = 16'h6180;
 buffer[276] = 16'h6147;
 buffer[277] = 16'h6147;
 buffer[278] = 16'h700C;
 buffer[279] = 16'h0220;
 buffer[280] = 16'h7242;
 buffer[281] = 16'h003E;
 buffer[282] = 16'h6B8D;
 buffer[283] = 16'h6B8D;
 buffer[284] = 16'h6180;
 buffer[285] = 16'h6147;
 buffer[286] = 16'h700C;
 buffer[287] = 16'h0230;
 buffer[288] = 16'h7242;
 buffer[289] = 16'h0040;
 buffer[290] = 16'h6B8D;
 buffer[291] = 16'h6B8D;
 buffer[292] = 16'h6081;
 buffer[293] = 16'h6147;
 buffer[294] = 16'h6180;
 buffer[295] = 16'h6147;
 buffer[296] = 16'h700C;
 buffer[297] = 16'h0240;
 buffer[298] = 16'h4001;
 buffer[299] = 16'h7C0C;
 buffer[300] = 16'h0254;
 buffer[301] = 16'h2101;
 buffer[302] = 16'h6023;
 buffer[303] = 16'h710F;
 buffer[304] = 16'h025A;
 buffer[305] = 16'h3C02;
 buffer[306] = 16'h003E;
 buffer[307] = 16'h721F;
 buffer[308] = 16'h0262;
 buffer[309] = 16'h3002;
 buffer[310] = 16'h003C;
 buffer[311] = 16'h781C;
 buffer[312] = 16'h026A;
 buffer[313] = 16'h3002;
 buffer[314] = 16'h003D;
 buffer[315] = 16'h701C;
 buffer[316] = 16'h0272;
 buffer[317] = 16'h3003;
 buffer[318] = 16'h3E3C;
 buffer[319] = 16'h711C;
 buffer[320] = 16'h027A;
 buffer[321] = 16'h3E01;
 buffer[322] = 16'h761F;
 buffer[323] = 16'h0282;
 buffer[324] = 16'h3002;
 buffer[325] = 16'h003E;
 buffer[326] = 16'h791C;
 buffer[327] = 16'h0288;
 buffer[328] = 16'h3E02;
 buffer[329] = 16'h003D;
 buffer[330] = 16'h7F1F;
 buffer[331] = 16'h0290;
 buffer[332] = 16'h7404;
 buffer[333] = 16'h6375;
 buffer[334] = 16'h006B;
 buffer[335] = 16'h6180;
 buffer[336] = 16'h718D;
 buffer[337] = 16'h0298;
 buffer[338] = 16'h2D04;
 buffer[339] = 16'h6F72;
 buffer[340] = 16'h0074;
 buffer[341] = 16'h6180;
 buffer[342] = 16'h6147;
 buffer[343] = 16'h6180;
 buffer[344] = 16'h6B8D;
 buffer[345] = 16'h700C;
 buffer[346] = 16'h02A4;
 buffer[347] = 16'h3202;
 buffer[348] = 16'h002F;
 buffer[349] = 16'h8001;
 buffer[350] = 16'h790F;
 buffer[351] = 16'h02B6;
 buffer[352] = 16'h3202;
 buffer[353] = 16'h002A;
 buffer[354] = 16'h741C;
 buffer[355] = 16'h02C0;
 buffer[356] = 16'h3102;
 buffer[357] = 16'h002B;
 buffer[358] = 16'h731C;
 buffer[359] = 16'h02C8;
 buffer[360] = 16'h7303;
 buffer[361] = 16'h4070;
 buffer[362] = 16'h6E81;
 buffer[363] = 16'h80FF;
 buffer[364] = 16'h730F;
 buffer[365] = 16'h02D0;
 buffer[366] = 16'h6507;
 buffer[367] = 16'h6578;
 buffer[368] = 16'h7563;
 buffer[369] = 16'h6574;
 buffer[370] = 16'h6147;
 buffer[371] = 16'h700C;
 buffer[372] = 16'h02DC;
 buffer[373] = 16'h6203;
 buffer[374] = 16'h6579;
 buffer[375] = 16'h8FFD;
 buffer[376] = 16'h6600;
 buffer[377] = 16'h6023;
 buffer[378] = 16'h710F;
 buffer[379] = 16'h02EA;
 buffer[380] = 16'h6302;
 buffer[381] = 16'h0040;
 buffer[382] = 16'h6081;
 buffer[383] = 16'h6C00;
 buffer[384] = 16'h6180;
 buffer[385] = 16'h8001;
 buffer[386] = 16'h6303;
 buffer[387] = 16'h2187;
 buffer[388] = 16'h8008;
 buffer[389] = 16'h6903;
 buffer[390] = 16'h0189;
 buffer[391] = 16'h80FF;
 buffer[392] = 16'h730F;
 buffer[393] = 16'h700C;
 buffer[394] = 16'h02F8;
 buffer[395] = 16'h6302;
 buffer[396] = 16'h0021;
 buffer[397] = 16'h6180;
 buffer[398] = 16'h80FF;
 buffer[399] = 16'h6303;
 buffer[400] = 16'h6081;
 buffer[401] = 16'h8008;
 buffer[402] = 16'h6D03;
 buffer[403] = 16'h6403;
 buffer[404] = 16'h6180;
 buffer[405] = 16'h414F;
 buffer[406] = 16'h6081;
 buffer[407] = 16'h6C00;
 buffer[408] = 16'h6180;
 buffer[409] = 16'h8001;
 buffer[410] = 16'h6303;
 buffer[411] = 16'h8000;
 buffer[412] = 16'h6703;
 buffer[413] = 16'h80FF;
 buffer[414] = 16'h6503;
 buffer[415] = 16'h6147;
 buffer[416] = 16'h6181;
 buffer[417] = 16'h6503;
 buffer[418] = 16'h6B8D;
 buffer[419] = 16'h6303;
 buffer[420] = 16'h6503;
 buffer[421] = 16'h6180;
 buffer[422] = 16'h6023;
 buffer[423] = 16'h710F;
 buffer[424] = 16'h0316;
 buffer[425] = 16'h7503;
 buffer[426] = 16'h2B6D;
 buffer[427] = 16'h6181;
 buffer[428] = 16'h6181;
 buffer[429] = 16'h6203;
 buffer[430] = 16'h6147;
 buffer[431] = 16'h6B81;
 buffer[432] = 16'h8000;
 buffer[433] = 16'h6F13;
 buffer[434] = 16'h6147;
 buffer[435] = 16'h6181;
 buffer[436] = 16'h6181;
 buffer[437] = 16'h6303;
 buffer[438] = 16'h6810;
 buffer[439] = 16'h6B8D;
 buffer[440] = 16'h6403;
 buffer[441] = 16'h6147;
 buffer[442] = 16'h6403;
 buffer[443] = 16'h6810;
 buffer[444] = 16'h6B8D;
 buffer[445] = 16'h6303;
 buffer[446] = 16'h6600;
 buffer[447] = 16'h6310;
 buffer[448] = 16'h6B8D;
 buffer[449] = 16'h718C;
 buffer[450] = 16'h0352;
 buffer[451] = 16'h6445;
 buffer[452] = 16'h766F;
 buffer[453] = 16'h7261;
 buffer[454] = 16'h6B8D;
 buffer[455] = 16'h700C;
 buffer[456] = 16'h0386;
 buffer[457] = 16'h7502;
 buffer[458] = 16'h0070;
 buffer[459] = 16'h41C6;
 buffer[460] = 16'h7E8C;
 buffer[461] = 16'h0392;
 buffer[462] = 16'h6446;
 buffer[463] = 16'h756F;
 buffer[464] = 16'h6573;
 buffer[465] = 16'h0072;
 buffer[466] = 16'h41CB;
 buffer[467] = 16'h6C00;
 buffer[468] = 16'h6B8D;
 buffer[469] = 16'h6C00;
 buffer[470] = 16'h720F;
 buffer[471] = 16'h039C;
 buffer[472] = 16'h6204;
 buffer[473] = 16'h7361;
 buffer[474] = 16'h0065;
 buffer[475] = 16'hFE80;
 buffer[476] = 16'h700C;
 buffer[477] = 16'h03B0;
 buffer[478] = 16'h7404;
 buffer[479] = 16'h6D65;
 buffer[480] = 16'h0070;
 buffer[481] = 16'hFE82;
 buffer[482] = 16'h700C;
 buffer[483] = 16'h03BC;
 buffer[484] = 16'h3E03;
 buffer[485] = 16'h6E69;
 buffer[486] = 16'hFE84;
 buffer[487] = 16'h700C;
 buffer[488] = 16'h03C8;
 buffer[489] = 16'h2304;
 buffer[490] = 16'h6974;
 buffer[491] = 16'h0062;
 buffer[492] = 16'hFE86;
 buffer[493] = 16'h700C;
 buffer[494] = 16'h03D2;
 buffer[495] = 16'h7403;
 buffer[496] = 16'h6269;
 buffer[497] = 16'hFE88;
 buffer[498] = 16'h700C;
 buffer[499] = 16'h03DE;
 buffer[500] = 16'h2705;
 buffer[501] = 16'h7665;
 buffer[502] = 16'h6C61;
 buffer[503] = 16'hFE8A;
 buffer[504] = 16'h700C;
 buffer[505] = 16'h03E8;
 buffer[506] = 16'h2706;
 buffer[507] = 16'h6261;
 buffer[508] = 16'h726F;
 buffer[509] = 16'h0074;
 buffer[510] = 16'hFE8C;
 buffer[511] = 16'h700C;
 buffer[512] = 16'h03F4;
 buffer[513] = 16'h6803;
 buffer[514] = 16'h646C;
 buffer[515] = 16'hFE8E;
 buffer[516] = 16'h700C;
 buffer[517] = 16'h0402;
 buffer[518] = 16'h6307;
 buffer[519] = 16'h6E6F;
 buffer[520] = 16'h6574;
 buffer[521] = 16'h7478;
 buffer[522] = 16'hFE90;
 buffer[523] = 16'h700C;
 buffer[524] = 16'h040C;
 buffer[525] = 16'h660E;
 buffer[526] = 16'h726F;
 buffer[527] = 16'h6874;
 buffer[528] = 16'h772D;
 buffer[529] = 16'h726F;
 buffer[530] = 16'h6C64;
 buffer[531] = 16'h7369;
 buffer[532] = 16'h0074;
 buffer[533] = 16'hFEA2;
 buffer[534] = 16'h700C;
 buffer[535] = 16'h041A;
 buffer[536] = 16'h6307;
 buffer[537] = 16'h7275;
 buffer[538] = 16'h6572;
 buffer[539] = 16'h746E;
 buffer[540] = 16'hFEA8;
 buffer[541] = 16'h700C;
 buffer[542] = 16'h0430;
 buffer[543] = 16'h6402;
 buffer[544] = 16'h0070;
 buffer[545] = 16'hFEAC;
 buffer[546] = 16'h700C;
 buffer[547] = 16'h043E;
 buffer[548] = 16'h6C04;
 buffer[549] = 16'h7361;
 buffer[550] = 16'h0074;
 buffer[551] = 16'hFEAE;
 buffer[552] = 16'h700C;
 buffer[553] = 16'h0448;
 buffer[554] = 16'h2705;
 buffer[555] = 16'h6B3F;
 buffer[556] = 16'h7965;
 buffer[557] = 16'hFEB0;
 buffer[558] = 16'h700C;
 buffer[559] = 16'h0454;
 buffer[560] = 16'h2705;
 buffer[561] = 16'h6D65;
 buffer[562] = 16'h7469;
 buffer[563] = 16'hFEB2;
 buffer[564] = 16'h700C;
 buffer[565] = 16'h0460;
 buffer[566] = 16'h2705;
 buffer[567] = 16'h6F62;
 buffer[568] = 16'h746F;
 buffer[569] = 16'hFEB4;
 buffer[570] = 16'h700C;
 buffer[571] = 16'h046C;
 buffer[572] = 16'h2702;
 buffer[573] = 16'h005C;
 buffer[574] = 16'hFEB6;
 buffer[575] = 16'h700C;
 buffer[576] = 16'h0478;
 buffer[577] = 16'h2706;
 buffer[578] = 16'h616E;
 buffer[579] = 16'h656D;
 buffer[580] = 16'h003F;
 buffer[581] = 16'hFEB8;
 buffer[582] = 16'h700C;
 buffer[583] = 16'h0482;
 buffer[584] = 16'h2704;
 buffer[585] = 16'h2C24;
 buffer[586] = 16'h006E;
 buffer[587] = 16'hFEBA;
 buffer[588] = 16'h700C;
 buffer[589] = 16'h0490;
 buffer[590] = 16'h2706;
 buffer[591] = 16'h766F;
 buffer[592] = 16'h7265;
 buffer[593] = 16'h0074;
 buffer[594] = 16'hFEBC;
 buffer[595] = 16'h700C;
 buffer[596] = 16'h049C;
 buffer[597] = 16'h2702;
 buffer[598] = 16'h003B;
 buffer[599] = 16'hFEBE;
 buffer[600] = 16'h700C;
 buffer[601] = 16'h04AA;
 buffer[602] = 16'h2707;
 buffer[603] = 16'h7263;
 buffer[604] = 16'h6165;
 buffer[605] = 16'h6574;
 buffer[606] = 16'hFEC0;
 buffer[607] = 16'h700C;
 buffer[608] = 16'h04B4;
 buffer[609] = 16'h3F04;
 buffer[610] = 16'h7564;
 buffer[611] = 16'h0070;
 buffer[612] = 16'h6081;
 buffer[613] = 16'h2267;
 buffer[614] = 16'h708D;
 buffer[615] = 16'h700C;
 buffer[616] = 16'h04C2;
 buffer[617] = 16'h7203;
 buffer[618] = 16'h746F;
 buffer[619] = 16'h6147;
 buffer[620] = 16'h6180;
 buffer[621] = 16'h6B8D;
 buffer[622] = 16'h718C;
 buffer[623] = 16'h04D2;
 buffer[624] = 16'h3205;
 buffer[625] = 16'h7264;
 buffer[626] = 16'h706F;
 buffer[627] = 16'h6103;
 buffer[628] = 16'h710F;
 buffer[629] = 16'h04E0;
 buffer[630] = 16'h3204;
 buffer[631] = 16'h7564;
 buffer[632] = 16'h0070;
 buffer[633] = 16'h6181;
 buffer[634] = 16'h718D;
 buffer[635] = 16'h04EC;
 buffer[636] = 16'h6E06;
 buffer[637] = 16'h6765;
 buffer[638] = 16'h7461;
 buffer[639] = 16'h0065;
 buffer[640] = 16'h7D1C;
 buffer[641] = 16'h04F8;
 buffer[642] = 16'h6407;
 buffer[643] = 16'h656E;
 buffer[644] = 16'h6167;
 buffer[645] = 16'h6574;
 buffer[646] = 16'h6600;
 buffer[647] = 16'h6147;
 buffer[648] = 16'h6600;
 buffer[649] = 16'h8001;
 buffer[650] = 16'h41AB;
 buffer[651] = 16'h6B8D;
 buffer[652] = 16'h720F;
 buffer[653] = 16'h0504;
 buffer[654] = 16'h2D01;
 buffer[655] = 16'h6D10;
 buffer[656] = 16'h720F;
 buffer[657] = 16'h051C;
 buffer[658] = 16'h6103;
 buffer[659] = 16'h7362;
 buffer[660] = 16'h7A1C;
 buffer[661] = 16'h0524;
 buffer[662] = 16'h6D03;
 buffer[663] = 16'h7861;
 buffer[664] = 16'h7B1F;
 buffer[665] = 16'h052C;
 buffer[666] = 16'h6D03;
 buffer[667] = 16'h6E69;
 buffer[668] = 16'h7C1F;
 buffer[669] = 16'h0534;
 buffer[670] = 16'h7706;
 buffer[671] = 16'h7469;
 buffer[672] = 16'h6968;
 buffer[673] = 16'h006E;
 buffer[674] = 16'h6181;
 buffer[675] = 16'h428F;
 buffer[676] = 16'h6147;
 buffer[677] = 16'h428F;
 buffer[678] = 16'h6B8D;
 buffer[679] = 16'h7F0F;
 buffer[680] = 16'h053C;
 buffer[681] = 16'h7506;
 buffer[682] = 16'h2F6D;
 buffer[683] = 16'h6F6D;
 buffer[684] = 16'h0064;
 buffer[685] = 16'h4279;
 buffer[686] = 16'h6F03;
 buffer[687] = 16'h22D6;
 buffer[688] = 16'h6D10;
 buffer[689] = 16'h800F;
 buffer[690] = 16'h6147;
 buffer[691] = 16'h6147;
 buffer[692] = 16'h6081;
 buffer[693] = 16'h41AB;
 buffer[694] = 16'h6147;
 buffer[695] = 16'h6147;
 buffer[696] = 16'h6081;
 buffer[697] = 16'h41AB;
 buffer[698] = 16'h6B8D;
 buffer[699] = 16'h6203;
 buffer[700] = 16'h6081;
 buffer[701] = 16'h6B8D;
 buffer[702] = 16'h6B81;
 buffer[703] = 16'h6180;
 buffer[704] = 16'h6147;
 buffer[705] = 16'h41AB;
 buffer[706] = 16'h6B8D;
 buffer[707] = 16'h6403;
 buffer[708] = 16'h22CA;
 buffer[709] = 16'h6147;
 buffer[710] = 16'h6103;
 buffer[711] = 16'h6310;
 buffer[712] = 16'h6B8D;
 buffer[713] = 16'h02CB;
 buffer[714] = 16'h6103;
 buffer[715] = 16'h6B8D;
 buffer[716] = 16'h6B81;
 buffer[717] = 16'h22D2;
 buffer[718] = 16'h6B8D;
 buffer[719] = 16'h6A00;
 buffer[720] = 16'h6147;
 buffer[721] = 16'h02B3;
 buffer[722] = 16'h6B8D;
 buffer[723] = 16'h6103;
 buffer[724] = 16'h6103;
 buffer[725] = 16'h718C;
 buffer[726] = 16'h6103;
 buffer[727] = 16'h4273;
 buffer[728] = 16'h8000;
 buffer[729] = 16'h6600;
 buffer[730] = 16'h708D;
 buffer[731] = 16'h0552;
 buffer[732] = 16'h6D05;
 buffer[733] = 16'h6D2F;
 buffer[734] = 16'h646F;
 buffer[735] = 16'h6081;
 buffer[736] = 16'h6810;
 buffer[737] = 16'h6081;
 buffer[738] = 16'h6147;
 buffer[739] = 16'h22E8;
 buffer[740] = 16'h6D10;
 buffer[741] = 16'h6147;
 buffer[742] = 16'h4286;
 buffer[743] = 16'h6B8D;
 buffer[744] = 16'h6147;
 buffer[745] = 16'h6081;
 buffer[746] = 16'h6810;
 buffer[747] = 16'h22EE;
 buffer[748] = 16'h6B81;
 buffer[749] = 16'h6203;
 buffer[750] = 16'h6B8D;
 buffer[751] = 16'h42AD;
 buffer[752] = 16'h6B8D;
 buffer[753] = 16'h22F5;
 buffer[754] = 16'h6180;
 buffer[755] = 16'h6D10;
 buffer[756] = 16'h718C;
 buffer[757] = 16'h700C;
 buffer[758] = 16'h05B8;
 buffer[759] = 16'h2F04;
 buffer[760] = 16'h6F6D;
 buffer[761] = 16'h0064;
 buffer[762] = 16'h6181;
 buffer[763] = 16'h6810;
 buffer[764] = 16'h6180;
 buffer[765] = 16'h02DF;
 buffer[766] = 16'h05EE;
 buffer[767] = 16'h6D03;
 buffer[768] = 16'h646F;
 buffer[769] = 16'h42FA;
 buffer[770] = 16'h710F;
 buffer[771] = 16'h05FE;
 buffer[772] = 16'h2F01;
 buffer[773] = 16'h42FA;
 buffer[774] = 16'h700F;
 buffer[775] = 16'h0608;
 buffer[776] = 16'h7503;
 buffer[777] = 16'h2A6D;
 buffer[778] = 16'h8000;
 buffer[779] = 16'h6180;
 buffer[780] = 16'h800F;
 buffer[781] = 16'h6147;
 buffer[782] = 16'h6081;
 buffer[783] = 16'h41AB;
 buffer[784] = 16'h6147;
 buffer[785] = 16'h6147;
 buffer[786] = 16'h6081;
 buffer[787] = 16'h41AB;
 buffer[788] = 16'h6B8D;
 buffer[789] = 16'h6203;
 buffer[790] = 16'h6B8D;
 buffer[791] = 16'h231D;
 buffer[792] = 16'h6147;
 buffer[793] = 16'h6181;
 buffer[794] = 16'h41AB;
 buffer[795] = 16'h6B8D;
 buffer[796] = 16'h6203;
 buffer[797] = 16'h6B81;
 buffer[798] = 16'h2323;
 buffer[799] = 16'h6B8D;
 buffer[800] = 16'h6A00;
 buffer[801] = 16'h6147;
 buffer[802] = 16'h030E;
 buffer[803] = 16'h6B8D;
 buffer[804] = 16'h6103;
 buffer[805] = 16'h426B;
 buffer[806] = 16'h710F;
 buffer[807] = 16'h0610;
 buffer[808] = 16'h2A01;
 buffer[809] = 16'h430A;
 buffer[810] = 16'h710F;
 buffer[811] = 16'h0650;
 buffer[812] = 16'h6D02;
 buffer[813] = 16'h002A;
 buffer[814] = 16'h4279;
 buffer[815] = 16'h6503;
 buffer[816] = 16'h6810;
 buffer[817] = 16'h6147;
 buffer[818] = 16'h6A10;
 buffer[819] = 16'h6180;
 buffer[820] = 16'h6A10;
 buffer[821] = 16'h430A;
 buffer[822] = 16'h6B8D;
 buffer[823] = 16'h2339;
 buffer[824] = 16'h0286;
 buffer[825] = 16'h700C;
 buffer[826] = 16'h0658;
 buffer[827] = 16'h2A05;
 buffer[828] = 16'h6D2F;
 buffer[829] = 16'h646F;
 buffer[830] = 16'h6147;
 buffer[831] = 16'h432E;
 buffer[832] = 16'h6B8D;
 buffer[833] = 16'h02DF;
 buffer[834] = 16'h0676;
 buffer[835] = 16'h2A02;
 buffer[836] = 16'h002F;
 buffer[837] = 16'h433E;
 buffer[838] = 16'h700F;
 buffer[839] = 16'h0686;
 buffer[840] = 16'h6305;
 buffer[841] = 16'h6C65;
 buffer[842] = 16'h2B6C;
 buffer[843] = 16'h8002;
 buffer[844] = 16'h720F;
 buffer[845] = 16'h0690;
 buffer[846] = 16'h6305;
 buffer[847] = 16'h6C65;
 buffer[848] = 16'h2D6C;
 buffer[849] = 16'h8002;
 buffer[850] = 16'h028F;
 buffer[851] = 16'h069C;
 buffer[852] = 16'h6305;
 buffer[853] = 16'h6C65;
 buffer[854] = 16'h736C;
 buffer[855] = 16'h8001;
 buffer[856] = 16'h7D0F;
 buffer[857] = 16'h06A8;
 buffer[858] = 16'h6202;
 buffer[859] = 16'h006C;
 buffer[860] = 16'h8020;
 buffer[861] = 16'h700C;
 buffer[862] = 16'h06B4;
 buffer[863] = 16'h3E05;
 buffer[864] = 16'h6863;
 buffer[865] = 16'h7261;
 buffer[866] = 16'h807F;
 buffer[867] = 16'h6303;
 buffer[868] = 16'h6081;
 buffer[869] = 16'h807F;
 buffer[870] = 16'h435C;
 buffer[871] = 16'h42A2;
 buffer[872] = 16'h236B;
 buffer[873] = 16'h6103;
 buffer[874] = 16'h805F;
 buffer[875] = 16'h700C;
 buffer[876] = 16'h700C;
 buffer[877] = 16'h06BE;
 buffer[878] = 16'h2B02;
 buffer[879] = 16'h0021;
 buffer[880] = 16'h414F;
 buffer[881] = 16'h6C00;
 buffer[882] = 16'h6203;
 buffer[883] = 16'h6180;
 buffer[884] = 16'h6023;
 buffer[885] = 16'h710F;
 buffer[886] = 16'h06DC;
 buffer[887] = 16'h3202;
 buffer[888] = 16'h0021;
 buffer[889] = 16'h6180;
 buffer[890] = 16'h6181;
 buffer[891] = 16'h6023;
 buffer[892] = 16'h6103;
 buffer[893] = 16'h434B;
 buffer[894] = 16'h6023;
 buffer[895] = 16'h710F;
 buffer[896] = 16'h06EE;
 buffer[897] = 16'h3202;
 buffer[898] = 16'h0040;
 buffer[899] = 16'h6081;
 buffer[900] = 16'h434B;
 buffer[901] = 16'h6C00;
 buffer[902] = 16'h6180;
 buffer[903] = 16'h7C0C;
 buffer[904] = 16'h0702;
 buffer[905] = 16'h6305;
 buffer[906] = 16'h756F;
 buffer[907] = 16'h746E;
 buffer[908] = 16'h6081;
 buffer[909] = 16'h6310;
 buffer[910] = 16'h6180;
 buffer[911] = 16'h017E;
 buffer[912] = 16'h0712;
 buffer[913] = 16'h6804;
 buffer[914] = 16'h7265;
 buffer[915] = 16'h0065;
 buffer[916] = 16'hFEAC;
 buffer[917] = 16'h7C0C;
 buffer[918] = 16'h0722;
 buffer[919] = 16'h6107;
 buffer[920] = 16'h696C;
 buffer[921] = 16'h6E67;
 buffer[922] = 16'h6465;
 buffer[923] = 16'h6081;
 buffer[924] = 16'h8000;
 buffer[925] = 16'h8002;
 buffer[926] = 16'h42AD;
 buffer[927] = 16'h6103;
 buffer[928] = 16'h6081;
 buffer[929] = 16'h23A5;
 buffer[930] = 16'h8002;
 buffer[931] = 16'h6180;
 buffer[932] = 16'h428F;
 buffer[933] = 16'h720F;
 buffer[934] = 16'h072E;
 buffer[935] = 16'h6105;
 buffer[936] = 16'h696C;
 buffer[937] = 16'h6E67;
 buffer[938] = 16'h4394;
 buffer[939] = 16'h439B;
 buffer[940] = 16'hFEAC;
 buffer[941] = 16'h6023;
 buffer[942] = 16'h710F;
 buffer[943] = 16'h074E;
 buffer[944] = 16'h7003;
 buffer[945] = 16'h6461;
 buffer[946] = 16'h4394;
 buffer[947] = 16'h8050;
 buffer[948] = 16'h6203;
 buffer[949] = 16'h039B;
 buffer[950] = 16'h0760;
 buffer[951] = 16'h4008;
 buffer[952] = 16'h7865;
 buffer[953] = 16'h6365;
 buffer[954] = 16'h7475;
 buffer[955] = 16'h0065;
 buffer[956] = 16'h6C00;
 buffer[957] = 16'h4264;
 buffer[958] = 16'h23C0;
 buffer[959] = 16'h0172;
 buffer[960] = 16'h700C;
 buffer[961] = 16'h076E;
 buffer[962] = 16'h6604;
 buffer[963] = 16'h6C69;
 buffer[964] = 16'h006C;
 buffer[965] = 16'h6180;
 buffer[966] = 16'h6147;
 buffer[967] = 16'h6180;
 buffer[968] = 16'h03CC;
 buffer[969] = 16'h4279;
 buffer[970] = 16'h418D;
 buffer[971] = 16'h6310;
 buffer[972] = 16'h6B81;
 buffer[973] = 16'h23D2;
 buffer[974] = 16'h6B8D;
 buffer[975] = 16'h6A00;
 buffer[976] = 16'h6147;
 buffer[977] = 16'h03C9;
 buffer[978] = 16'h6B8D;
 buffer[979] = 16'h6103;
 buffer[980] = 16'h0273;
 buffer[981] = 16'h0784;
 buffer[982] = 16'h6505;
 buffer[983] = 16'h6172;
 buffer[984] = 16'h6573;
 buffer[985] = 16'h8000;
 buffer[986] = 16'h03C5;
 buffer[987] = 16'h07AC;
 buffer[988] = 16'h6405;
 buffer[989] = 16'h6769;
 buffer[990] = 16'h7469;
 buffer[991] = 16'h8009;
 buffer[992] = 16'h6181;
 buffer[993] = 16'h6803;
 buffer[994] = 16'h8007;
 buffer[995] = 16'h6303;
 buffer[996] = 16'h6203;
 buffer[997] = 16'h8030;
 buffer[998] = 16'h720F;
 buffer[999] = 16'h07B8;
 buffer[1000] = 16'h6507;
 buffer[1001] = 16'h7478;
 buffer[1002] = 16'h6172;
 buffer[1003] = 16'h7463;
 buffer[1004] = 16'h8000;
 buffer[1005] = 16'h6180;
 buffer[1006] = 16'h42AD;
 buffer[1007] = 16'h6180;
 buffer[1008] = 16'h03DF;
 buffer[1009] = 16'h07D0;
 buffer[1010] = 16'h3C02;
 buffer[1011] = 16'h0023;
 buffer[1012] = 16'h43B2;
 buffer[1013] = 16'hFE8E;
 buffer[1014] = 16'h6023;
 buffer[1015] = 16'h710F;
 buffer[1016] = 16'h07E4;
 buffer[1017] = 16'h6804;
 buffer[1018] = 16'h6C6F;
 buffer[1019] = 16'h0064;
 buffer[1020] = 16'hFE8E;
 buffer[1021] = 16'h6C00;
 buffer[1022] = 16'h6A00;
 buffer[1023] = 16'h6081;
 buffer[1024] = 16'hFE8E;
 buffer[1025] = 16'h6023;
 buffer[1026] = 16'h6103;
 buffer[1027] = 16'h018D;
 buffer[1028] = 16'h07F2;
 buffer[1029] = 16'h2301;
 buffer[1030] = 16'hFE80;
 buffer[1031] = 16'h6C00;
 buffer[1032] = 16'h43EC;
 buffer[1033] = 16'h03FC;
 buffer[1034] = 16'h080A;
 buffer[1035] = 16'h2302;
 buffer[1036] = 16'h0073;
 buffer[1037] = 16'h4406;
 buffer[1038] = 16'h6081;
 buffer[1039] = 16'h2411;
 buffer[1040] = 16'h040D;
 buffer[1041] = 16'h700C;
 buffer[1042] = 16'h0816;
 buffer[1043] = 16'h7304;
 buffer[1044] = 16'h6769;
 buffer[1045] = 16'h006E;
 buffer[1046] = 16'h6810;
 buffer[1047] = 16'h241A;
 buffer[1048] = 16'h802D;
 buffer[1049] = 16'h03FC;
 buffer[1050] = 16'h700C;
 buffer[1051] = 16'h0826;
 buffer[1052] = 16'h2302;
 buffer[1053] = 16'h003E;
 buffer[1054] = 16'h6103;
 buffer[1055] = 16'hFE8E;
 buffer[1056] = 16'h6C00;
 buffer[1057] = 16'h43B2;
 buffer[1058] = 16'h6181;
 buffer[1059] = 16'h028F;
 buffer[1060] = 16'h0838;
 buffer[1061] = 16'h7303;
 buffer[1062] = 16'h7274;
 buffer[1063] = 16'h6081;
 buffer[1064] = 16'h6147;
 buffer[1065] = 16'h6A10;
 buffer[1066] = 16'h43F4;
 buffer[1067] = 16'h440D;
 buffer[1068] = 16'h6B8D;
 buffer[1069] = 16'h4416;
 buffer[1070] = 16'h041E;
 buffer[1071] = 16'h084A;
 buffer[1072] = 16'h6803;
 buffer[1073] = 16'h7865;
 buffer[1074] = 16'h8010;
 buffer[1075] = 16'hFE80;
 buffer[1076] = 16'h6023;
 buffer[1077] = 16'h710F;
 buffer[1078] = 16'h0860;
 buffer[1079] = 16'h6407;
 buffer[1080] = 16'h6365;
 buffer[1081] = 16'h6D69;
 buffer[1082] = 16'h6C61;
 buffer[1083] = 16'h800A;
 buffer[1084] = 16'hFE80;
 buffer[1085] = 16'h6023;
 buffer[1086] = 16'h710F;
 buffer[1087] = 16'h086E;
 buffer[1088] = 16'h6406;
 buffer[1089] = 16'h6769;
 buffer[1090] = 16'h7469;
 buffer[1091] = 16'h003F;
 buffer[1092] = 16'h6147;
 buffer[1093] = 16'h8030;
 buffer[1094] = 16'h428F;
 buffer[1095] = 16'h8009;
 buffer[1096] = 16'h6181;
 buffer[1097] = 16'h6803;
 buffer[1098] = 16'h2457;
 buffer[1099] = 16'h6081;
 buffer[1100] = 16'h8020;
 buffer[1101] = 16'h6613;
 buffer[1102] = 16'h2451;
 buffer[1103] = 16'h8020;
 buffer[1104] = 16'h428F;
 buffer[1105] = 16'h8007;
 buffer[1106] = 16'h428F;
 buffer[1107] = 16'h6081;
 buffer[1108] = 16'h800A;
 buffer[1109] = 16'h6803;
 buffer[1110] = 16'h6403;
 buffer[1111] = 16'h6081;
 buffer[1112] = 16'h6B8D;
 buffer[1113] = 16'h7F0F;
 buffer[1114] = 16'h0880;
 buffer[1115] = 16'h6E07;
 buffer[1116] = 16'h6D75;
 buffer[1117] = 16'h6562;
 buffer[1118] = 16'h3F72;
 buffer[1119] = 16'hFE80;
 buffer[1120] = 16'h6C00;
 buffer[1121] = 16'h6147;
 buffer[1122] = 16'h8000;
 buffer[1123] = 16'h6181;
 buffer[1124] = 16'h438C;
 buffer[1125] = 16'h6181;
 buffer[1126] = 16'h417E;
 buffer[1127] = 16'h8024;
 buffer[1128] = 16'h6703;
 buffer[1129] = 16'h246F;
 buffer[1130] = 16'h4432;
 buffer[1131] = 16'h6180;
 buffer[1132] = 16'h6310;
 buffer[1133] = 16'h6180;
 buffer[1134] = 16'h6A00;
 buffer[1135] = 16'h6181;
 buffer[1136] = 16'h417E;
 buffer[1137] = 16'h802D;
 buffer[1138] = 16'h6703;
 buffer[1139] = 16'h6147;
 buffer[1140] = 16'h6180;
 buffer[1141] = 16'h6B81;
 buffer[1142] = 16'h428F;
 buffer[1143] = 16'h6180;
 buffer[1144] = 16'h6B81;
 buffer[1145] = 16'h6203;
 buffer[1146] = 16'h4264;
 buffer[1147] = 16'h24A0;
 buffer[1148] = 16'h6A00;
 buffer[1149] = 16'h6147;
 buffer[1150] = 16'h6081;
 buffer[1151] = 16'h6147;
 buffer[1152] = 16'h417E;
 buffer[1153] = 16'hFE80;
 buffer[1154] = 16'h6C00;
 buffer[1155] = 16'h4444;
 buffer[1156] = 16'h249A;
 buffer[1157] = 16'h6180;
 buffer[1158] = 16'hFE80;
 buffer[1159] = 16'h6C00;
 buffer[1160] = 16'h4329;
 buffer[1161] = 16'h6203;
 buffer[1162] = 16'h6B8D;
 buffer[1163] = 16'h6310;
 buffer[1164] = 16'h6B81;
 buffer[1165] = 16'h2492;
 buffer[1166] = 16'h6B8D;
 buffer[1167] = 16'h6A00;
 buffer[1168] = 16'h6147;
 buffer[1169] = 16'h047E;
 buffer[1170] = 16'h6B8D;
 buffer[1171] = 16'h6103;
 buffer[1172] = 16'h6B81;
 buffer[1173] = 16'h6003;
 buffer[1174] = 16'h2498;
 buffer[1175] = 16'h6D10;
 buffer[1176] = 16'h6180;
 buffer[1177] = 16'h049F;
 buffer[1178] = 16'h6B8D;
 buffer[1179] = 16'h6B8D;
 buffer[1180] = 16'h4273;
 buffer[1181] = 16'h4273;
 buffer[1182] = 16'h8000;
 buffer[1183] = 16'h6081;
 buffer[1184] = 16'h6B8D;
 buffer[1185] = 16'h4273;
 buffer[1186] = 16'h6B8D;
 buffer[1187] = 16'hFE80;
 buffer[1188] = 16'h6023;
 buffer[1189] = 16'h710F;
 buffer[1190] = 16'h08B6;
 buffer[1191] = 16'h3F03;
 buffer[1192] = 16'h7872;
 buffer[1193] = 16'h8FFE;
 buffer[1194] = 16'h6600;
 buffer[1195] = 16'h6C00;
 buffer[1196] = 16'h8001;
 buffer[1197] = 16'h6303;
 buffer[1198] = 16'h711C;
 buffer[1199] = 16'h094E;
 buffer[1200] = 16'h7403;
 buffer[1201] = 16'h2178;
 buffer[1202] = 16'h8FFE;
 buffer[1203] = 16'h6600;
 buffer[1204] = 16'h6C00;
 buffer[1205] = 16'h8002;
 buffer[1206] = 16'h6303;
 buffer[1207] = 16'h6010;
 buffer[1208] = 16'h24B2;
 buffer[1209] = 16'h8FFF;
 buffer[1210] = 16'h6600;
 buffer[1211] = 16'h6023;
 buffer[1212] = 16'h710F;
 buffer[1213] = 16'h0960;
 buffer[1214] = 16'h3F04;
 buffer[1215] = 16'h656B;
 buffer[1216] = 16'h0079;
 buffer[1217] = 16'hFEB0;
 buffer[1218] = 16'h03BC;
 buffer[1219] = 16'h097C;
 buffer[1220] = 16'h6504;
 buffer[1221] = 16'h696D;
 buffer[1222] = 16'h0074;
 buffer[1223] = 16'hFEB2;
 buffer[1224] = 16'h03BC;
 buffer[1225] = 16'h0988;
 buffer[1226] = 16'h6B03;
 buffer[1227] = 16'h7965;
 buffer[1228] = 16'h44C1;
 buffer[1229] = 16'h24CC;
 buffer[1230] = 16'h8FFF;
 buffer[1231] = 16'h6600;
 buffer[1232] = 16'h7C0C;
 buffer[1233] = 16'h0994;
 buffer[1234] = 16'h6E04;
 buffer[1235] = 16'h6675;
 buffer[1236] = 16'h003F;
 buffer[1237] = 16'h44C1;
 buffer[1238] = 16'h6081;
 buffer[1239] = 16'h24DC;
 buffer[1240] = 16'h6103;
 buffer[1241] = 16'h44CC;
 buffer[1242] = 16'h800D;
 buffer[1243] = 16'h770F;
 buffer[1244] = 16'h700C;
 buffer[1245] = 16'h09A4;
 buffer[1246] = 16'h7406;
 buffer[1247] = 16'h6D69;
 buffer[1248] = 16'h7265;
 buffer[1249] = 16'h0040;
 buffer[1250] = 16'h8FFB;
 buffer[1251] = 16'h6600;
 buffer[1252] = 16'h7C0C;
 buffer[1253] = 16'h09BC;
 buffer[1254] = 16'h7204;
 buffer[1255] = 16'h6267;
 buffer[1256] = 16'h0040;
 buffer[1257] = 16'h8FFD;
 buffer[1258] = 16'h6600;
 buffer[1259] = 16'h7C0C;
 buffer[1260] = 16'h09CC;
 buffer[1261] = 16'h7204;
 buffer[1262] = 16'h6267;
 buffer[1263] = 16'h0021;
 buffer[1264] = 16'h8FFD;
 buffer[1265] = 16'h6600;
 buffer[1266] = 16'h6023;
 buffer[1267] = 16'h710F;
 buffer[1268] = 16'h09DA;
 buffer[1269] = 16'h6208;
 buffer[1270] = 16'h7475;
 buffer[1271] = 16'h6F74;
 buffer[1272] = 16'h736E;
 buffer[1273] = 16'h0040;
 buffer[1274] = 16'h8FFC;
 buffer[1275] = 16'h6600;
 buffer[1276] = 16'h7C0C;
 buffer[1277] = 16'h09EA;
 buffer[1278] = 16'h7305;
 buffer[1279] = 16'h6170;
 buffer[1280] = 16'h6563;
 buffer[1281] = 16'h435C;
 buffer[1282] = 16'h04C7;
 buffer[1283] = 16'h09FC;
 buffer[1284] = 16'h7306;
 buffer[1285] = 16'h6170;
 buffer[1286] = 16'h6563;
 buffer[1287] = 16'h0073;
 buffer[1288] = 16'h8000;
 buffer[1289] = 16'h6B13;
 buffer[1290] = 16'h6147;
 buffer[1291] = 16'h050D;
 buffer[1292] = 16'h4501;
 buffer[1293] = 16'h6B81;
 buffer[1294] = 16'h2513;
 buffer[1295] = 16'h6B8D;
 buffer[1296] = 16'h6A00;
 buffer[1297] = 16'h6147;
 buffer[1298] = 16'h050C;
 buffer[1299] = 16'h6B8D;
 buffer[1300] = 16'h710F;
 buffer[1301] = 16'h0A08;
 buffer[1302] = 16'h7404;
 buffer[1303] = 16'h7079;
 buffer[1304] = 16'h0065;
 buffer[1305] = 16'h6147;
 buffer[1306] = 16'h051D;
 buffer[1307] = 16'h438C;
 buffer[1308] = 16'h44C7;
 buffer[1309] = 16'h6B81;
 buffer[1310] = 16'h2523;
 buffer[1311] = 16'h6B8D;
 buffer[1312] = 16'h6A00;
 buffer[1313] = 16'h6147;
 buffer[1314] = 16'h051B;
 buffer[1315] = 16'h6B8D;
 buffer[1316] = 16'h6103;
 buffer[1317] = 16'h710F;
 buffer[1318] = 16'h0A2C;
 buffer[1319] = 16'h6302;
 buffer[1320] = 16'h0072;
 buffer[1321] = 16'h800D;
 buffer[1322] = 16'h44C7;
 buffer[1323] = 16'h800A;
 buffer[1324] = 16'h04C7;
 buffer[1325] = 16'h0A4E;
 buffer[1326] = 16'h6443;
 buffer[1327] = 16'h246F;
 buffer[1328] = 16'h6B8D;
 buffer[1329] = 16'h6B81;
 buffer[1330] = 16'h6B8D;
 buffer[1331] = 16'h438C;
 buffer[1332] = 16'h6203;
 buffer[1333] = 16'h439B;
 buffer[1334] = 16'h6147;
 buffer[1335] = 16'h6180;
 buffer[1336] = 16'h6147;
 buffer[1337] = 16'h700C;
 buffer[1338] = 16'h0A5C;
 buffer[1339] = 16'h2443;
 buffer[1340] = 16'h7C22;
 buffer[1341] = 16'h4530;
 buffer[1342] = 16'h700C;
 buffer[1343] = 16'h0A76;
 buffer[1344] = 16'h2E02;
 buffer[1345] = 16'h0024;
 buffer[1346] = 16'h438C;
 buffer[1347] = 16'h0519;
 buffer[1348] = 16'h0A80;
 buffer[1349] = 16'h2E43;
 buffer[1350] = 16'h7C22;
 buffer[1351] = 16'h4530;
 buffer[1352] = 16'h0542;
 buffer[1353] = 16'h0A8A;
 buffer[1354] = 16'h2E02;
 buffer[1355] = 16'h0072;
 buffer[1356] = 16'h6147;
 buffer[1357] = 16'h4427;
 buffer[1358] = 16'h6B8D;
 buffer[1359] = 16'h6181;
 buffer[1360] = 16'h428F;
 buffer[1361] = 16'h4508;
 buffer[1362] = 16'h0519;
 buffer[1363] = 16'h0A94;
 buffer[1364] = 16'h7503;
 buffer[1365] = 16'h722E;
 buffer[1366] = 16'h6147;
 buffer[1367] = 16'h43F4;
 buffer[1368] = 16'h440D;
 buffer[1369] = 16'h441E;
 buffer[1370] = 16'h6B8D;
 buffer[1371] = 16'h6181;
 buffer[1372] = 16'h428F;
 buffer[1373] = 16'h4508;
 buffer[1374] = 16'h0519;
 buffer[1375] = 16'h0AA8;
 buffer[1376] = 16'h7502;
 buffer[1377] = 16'h002E;
 buffer[1378] = 16'h43F4;
 buffer[1379] = 16'h440D;
 buffer[1380] = 16'h441E;
 buffer[1381] = 16'h4501;
 buffer[1382] = 16'h0519;
 buffer[1383] = 16'h0AC0;
 buffer[1384] = 16'h2E01;
 buffer[1385] = 16'hFE80;
 buffer[1386] = 16'h6C00;
 buffer[1387] = 16'h800A;
 buffer[1388] = 16'h6503;
 buffer[1389] = 16'h256F;
 buffer[1390] = 16'h0562;
 buffer[1391] = 16'h4427;
 buffer[1392] = 16'h4501;
 buffer[1393] = 16'h0519;
 buffer[1394] = 16'h0AD0;
 buffer[1395] = 16'h2E02;
 buffer[1396] = 16'h0023;
 buffer[1397] = 16'hFE80;
 buffer[1398] = 16'h6C00;
 buffer[1399] = 16'h6180;
 buffer[1400] = 16'h443B;
 buffer[1401] = 16'h4569;
 buffer[1402] = 16'hFE80;
 buffer[1403] = 16'h6023;
 buffer[1404] = 16'h710F;
 buffer[1405] = 16'h0AE6;
 buffer[1406] = 16'h7503;
 buffer[1407] = 16'h232E;
 buffer[1408] = 16'hFE80;
 buffer[1409] = 16'h6C00;
 buffer[1410] = 16'h6180;
 buffer[1411] = 16'h443B;
 buffer[1412] = 16'h43F4;
 buffer[1413] = 16'h440D;
 buffer[1414] = 16'h441E;
 buffer[1415] = 16'h4501;
 buffer[1416] = 16'h4519;
 buffer[1417] = 16'hFE80;
 buffer[1418] = 16'h6023;
 buffer[1419] = 16'h710F;
 buffer[1420] = 16'h0AFC;
 buffer[1421] = 16'h7504;
 buffer[1422] = 16'h722E;
 buffer[1423] = 16'h0023;
 buffer[1424] = 16'hFE80;
 buffer[1425] = 16'h6C00;
 buffer[1426] = 16'h426B;
 buffer[1427] = 16'h426B;
 buffer[1428] = 16'h443B;
 buffer[1429] = 16'h6147;
 buffer[1430] = 16'h43F4;
 buffer[1431] = 16'h440D;
 buffer[1432] = 16'h441E;
 buffer[1433] = 16'h6B8D;
 buffer[1434] = 16'h6181;
 buffer[1435] = 16'h428F;
 buffer[1436] = 16'h4508;
 buffer[1437] = 16'h4519;
 buffer[1438] = 16'hFE80;
 buffer[1439] = 16'h6023;
 buffer[1440] = 16'h710F;
 buffer[1441] = 16'h0B1A;
 buffer[1442] = 16'h2E03;
 buffer[1443] = 16'h2372;
 buffer[1444] = 16'hFE80;
 buffer[1445] = 16'h6C00;
 buffer[1446] = 16'h426B;
 buffer[1447] = 16'h426B;
 buffer[1448] = 16'h443B;
 buffer[1449] = 16'h6147;
 buffer[1450] = 16'h4427;
 buffer[1451] = 16'h6B8D;
 buffer[1452] = 16'h6181;
 buffer[1453] = 16'h428F;
 buffer[1454] = 16'h4508;
 buffer[1455] = 16'h4519;
 buffer[1456] = 16'hFE80;
 buffer[1457] = 16'h6023;
 buffer[1458] = 16'h710F;
 buffer[1459] = 16'h0B44;
 buffer[1460] = 16'h6305;
 buffer[1461] = 16'h6F6D;
 buffer[1462] = 16'h6576;
 buffer[1463] = 16'h6147;
 buffer[1464] = 16'h05C1;
 buffer[1465] = 16'h6147;
 buffer[1466] = 16'h6081;
 buffer[1467] = 16'h417E;
 buffer[1468] = 16'h6B81;
 buffer[1469] = 16'h418D;
 buffer[1470] = 16'h6310;
 buffer[1471] = 16'h6B8D;
 buffer[1472] = 16'h6310;
 buffer[1473] = 16'h6B81;
 buffer[1474] = 16'h25C7;
 buffer[1475] = 16'h6B8D;
 buffer[1476] = 16'h6A00;
 buffer[1477] = 16'h6147;
 buffer[1478] = 16'h05B9;
 buffer[1479] = 16'h6B8D;
 buffer[1480] = 16'h6103;
 buffer[1481] = 16'h0273;
 buffer[1482] = 16'h0B68;
 buffer[1483] = 16'h7005;
 buffer[1484] = 16'h6361;
 buffer[1485] = 16'h246B;
 buffer[1486] = 16'h6081;
 buffer[1487] = 16'h6147;
 buffer[1488] = 16'h4279;
 buffer[1489] = 16'h6023;
 buffer[1490] = 16'h6103;
 buffer[1491] = 16'h6310;
 buffer[1492] = 16'h6180;
 buffer[1493] = 16'h45B7;
 buffer[1494] = 16'h6B8D;
 buffer[1495] = 16'h700C;
 buffer[1496] = 16'h0B96;
 buffer[1497] = 16'h3F01;
 buffer[1498] = 16'h6C00;
 buffer[1499] = 16'h0569;
 buffer[1500] = 16'h0BB2;
 buffer[1501] = 16'h3205;
 buffer[1502] = 16'h766F;
 buffer[1503] = 16'h7265;
 buffer[1504] = 16'h6147;
 buffer[1505] = 16'h6147;
 buffer[1506] = 16'h4279;
 buffer[1507] = 16'h6B8D;
 buffer[1508] = 16'h6B8D;
 buffer[1509] = 16'h426B;
 buffer[1510] = 16'h6147;
 buffer[1511] = 16'h426B;
 buffer[1512] = 16'h6B8D;
 buffer[1513] = 16'h700C;
 buffer[1514] = 16'h0BBA;
 buffer[1515] = 16'h3205;
 buffer[1516] = 16'h7773;
 buffer[1517] = 16'h7061;
 buffer[1518] = 16'h426B;
 buffer[1519] = 16'h6147;
 buffer[1520] = 16'h426B;
 buffer[1521] = 16'h6B8D;
 buffer[1522] = 16'h700C;
 buffer[1523] = 16'h0BD6;
 buffer[1524] = 16'h3204;
 buffer[1525] = 16'h696E;
 buffer[1526] = 16'h0070;
 buffer[1527] = 16'h426B;
 buffer[1528] = 16'h6103;
 buffer[1529] = 16'h426B;
 buffer[1530] = 16'h710F;
 buffer[1531] = 16'h0BE8;
 buffer[1532] = 16'h3204;
 buffer[1533] = 16'h6F72;
 buffer[1534] = 16'h0074;
 buffer[1535] = 16'h6180;
 buffer[1536] = 16'h6147;
 buffer[1537] = 16'h6147;
 buffer[1538] = 16'h45EE;
 buffer[1539] = 16'h6B8D;
 buffer[1540] = 16'h6B8D;
 buffer[1541] = 16'h6180;
 buffer[1542] = 16'h05EE;
 buffer[1543] = 16'h0BF8;
 buffer[1544] = 16'h6402;
 buffer[1545] = 16'h003D;
 buffer[1546] = 16'h6147;
 buffer[1547] = 16'h426B;
 buffer[1548] = 16'h6503;
 buffer[1549] = 16'h6180;
 buffer[1550] = 16'h6B8D;
 buffer[1551] = 16'h6503;
 buffer[1552] = 16'h6403;
 buffer[1553] = 16'h701C;
 buffer[1554] = 16'h0C10;
 buffer[1555] = 16'h6403;
 buffer[1556] = 16'h3E3C;
 buffer[1557] = 16'h460A;
 buffer[1558] = 16'h760C;
 buffer[1559] = 16'h0C26;
 buffer[1560] = 16'h6402;
 buffer[1561] = 16'h002B;
 buffer[1562] = 16'h426B;
 buffer[1563] = 16'h6203;
 buffer[1564] = 16'h6147;
 buffer[1565] = 16'h6181;
 buffer[1566] = 16'h6203;
 buffer[1567] = 16'h6081;
 buffer[1568] = 16'h426B;
 buffer[1569] = 16'h6F03;
 buffer[1570] = 16'h2626;
 buffer[1571] = 16'h6B8D;
 buffer[1572] = 16'h6310;
 buffer[1573] = 16'h0627;
 buffer[1574] = 16'h6B8D;
 buffer[1575] = 16'h700C;
 buffer[1576] = 16'h0C30;
 buffer[1577] = 16'h6402;
 buffer[1578] = 16'h002D;
 buffer[1579] = 16'h4286;
 buffer[1580] = 16'h061A;
 buffer[1581] = 16'h0C52;
 buffer[1582] = 16'h7303;
 buffer[1583] = 16'h643E;
 buffer[1584] = 16'h6081;
 buffer[1585] = 16'h781C;
 buffer[1586] = 16'h0C5C;
 buffer[1587] = 16'h6403;
 buffer[1588] = 16'h2B31;
 buffer[1589] = 16'h8001;
 buffer[1590] = 16'h4630;
 buffer[1591] = 16'h061A;
 buffer[1592] = 16'h0C66;
 buffer[1593] = 16'h6404;
 buffer[1594] = 16'h6F78;
 buffer[1595] = 16'h0072;
 buffer[1596] = 16'h426B;
 buffer[1597] = 16'h6503;
 buffer[1598] = 16'h4155;
 buffer[1599] = 16'h6503;
 buffer[1600] = 16'h718C;
 buffer[1601] = 16'h0C72;
 buffer[1602] = 16'h6404;
 buffer[1603] = 16'h6E61;
 buffer[1604] = 16'h0064;
 buffer[1605] = 16'h426B;
 buffer[1606] = 16'h6303;
 buffer[1607] = 16'h4155;
 buffer[1608] = 16'h6303;
 buffer[1609] = 16'h718C;
 buffer[1610] = 16'h0C84;
 buffer[1611] = 16'h6403;
 buffer[1612] = 16'h726F;
 buffer[1613] = 16'h426B;
 buffer[1614] = 16'h6403;
 buffer[1615] = 16'h4155;
 buffer[1616] = 16'h6403;
 buffer[1617] = 16'h718C;
 buffer[1618] = 16'h0C96;
 buffer[1619] = 16'h6407;
 buffer[1620] = 16'h6E69;
 buffer[1621] = 16'h6576;
 buffer[1622] = 16'h7472;
 buffer[1623] = 16'h6600;
 buffer[1624] = 16'h6180;
 buffer[1625] = 16'h6600;
 buffer[1626] = 16'h718C;
 buffer[1627] = 16'h0CA6;
 buffer[1628] = 16'h6402;
 buffer[1629] = 16'h003C;
 buffer[1630] = 16'h426B;
 buffer[1631] = 16'h4279;
 buffer[1632] = 16'h6703;
 buffer[1633] = 16'h2665;
 buffer[1634] = 16'h4273;
 buffer[1635] = 16'h6F03;
 buffer[1636] = 16'h0667;
 buffer[1637] = 16'h45F7;
 buffer[1638] = 16'h761F;
 buffer[1639] = 16'h0CB8;
 buffer[1640] = 16'h6402;
 buffer[1641] = 16'h003E;
 buffer[1642] = 16'h45EE;
 buffer[1643] = 16'h065E;
 buffer[1644] = 16'h0CD0;
 buffer[1645] = 16'h6403;
 buffer[1646] = 16'h3D30;
 buffer[1647] = 16'h6403;
 buffer[1648] = 16'h701C;
 buffer[1649] = 16'h0CDA;
 buffer[1650] = 16'h6403;
 buffer[1651] = 16'h3C30;
 buffer[1652] = 16'h8000;
 buffer[1653] = 16'h4630;
 buffer[1654] = 16'h065E;
 buffer[1655] = 16'h0CE4;
 buffer[1656] = 16'h6404;
 buffer[1657] = 16'h3C30;
 buffer[1658] = 16'h003E;
 buffer[1659] = 16'h466F;
 buffer[1660] = 16'h760C;
 buffer[1661] = 16'h0CF0;
 buffer[1662] = 16'h6403;
 buffer[1663] = 16'h2A32;
 buffer[1664] = 16'h4279;
 buffer[1665] = 16'h061A;
 buffer[1666] = 16'h0CFC;
 buffer[1667] = 16'h6403;
 buffer[1668] = 16'h2F32;
 buffer[1669] = 16'h6081;
 buffer[1670] = 16'h800F;
 buffer[1671] = 16'h6D03;
 buffer[1672] = 16'h6147;
 buffer[1673] = 16'h415D;
 buffer[1674] = 16'h6180;
 buffer[1675] = 16'h415D;
 buffer[1676] = 16'h6B8D;
 buffer[1677] = 16'h6403;
 buffer[1678] = 16'h718C;
 buffer[1679] = 16'h0D06;
 buffer[1680] = 16'h6403;
 buffer[1681] = 16'h2D31;
 buffer[1682] = 16'h8001;
 buffer[1683] = 16'h4630;
 buffer[1684] = 16'h4286;
 buffer[1685] = 16'h061A;
 buffer[1686] = 16'h0D20;
 buffer[1687] = 16'h2807;
 buffer[1688] = 16'h6170;
 buffer[1689] = 16'h7372;
 buffer[1690] = 16'h2965;
 buffer[1691] = 16'hFE82;
 buffer[1692] = 16'h6023;
 buffer[1693] = 16'h6103;
 buffer[1694] = 16'h6181;
 buffer[1695] = 16'h6147;
 buffer[1696] = 16'h6081;
 buffer[1697] = 16'h26E6;
 buffer[1698] = 16'h6A00;
 buffer[1699] = 16'hFE82;
 buffer[1700] = 16'h6C00;
 buffer[1701] = 16'h435C;
 buffer[1702] = 16'h6703;
 buffer[1703] = 16'h26C2;
 buffer[1704] = 16'h6147;
 buffer[1705] = 16'h438C;
 buffer[1706] = 16'hFE82;
 buffer[1707] = 16'h6C00;
 buffer[1708] = 16'h6180;
 buffer[1709] = 16'h428F;
 buffer[1710] = 16'h6810;
 buffer[1711] = 16'h6600;
 buffer[1712] = 16'h6B81;
 buffer[1713] = 16'h6910;
 buffer[1714] = 16'h6303;
 buffer[1715] = 16'h26C0;
 buffer[1716] = 16'h6B81;
 buffer[1717] = 16'h26BA;
 buffer[1718] = 16'h6B8D;
 buffer[1719] = 16'h6A00;
 buffer[1720] = 16'h6147;
 buffer[1721] = 16'h06A9;
 buffer[1722] = 16'h6B8D;
 buffer[1723] = 16'h6103;
 buffer[1724] = 16'h6B8D;
 buffer[1725] = 16'h6103;
 buffer[1726] = 16'h8000;
 buffer[1727] = 16'h708D;
 buffer[1728] = 16'h6A00;
 buffer[1729] = 16'h6B8D;
 buffer[1730] = 16'h6181;
 buffer[1731] = 16'h6180;
 buffer[1732] = 16'h6147;
 buffer[1733] = 16'h438C;
 buffer[1734] = 16'hFE82;
 buffer[1735] = 16'h6C00;
 buffer[1736] = 16'h6180;
 buffer[1737] = 16'h428F;
 buffer[1738] = 16'hFE82;
 buffer[1739] = 16'h6C00;
 buffer[1740] = 16'h435C;
 buffer[1741] = 16'h6703;
 buffer[1742] = 16'h26D0;
 buffer[1743] = 16'h6810;
 buffer[1744] = 16'h26DC;
 buffer[1745] = 16'h6B81;
 buffer[1746] = 16'h26D7;
 buffer[1747] = 16'h6B8D;
 buffer[1748] = 16'h6A00;
 buffer[1749] = 16'h6147;
 buffer[1750] = 16'h06C5;
 buffer[1751] = 16'h6B8D;
 buffer[1752] = 16'h6103;
 buffer[1753] = 16'h6081;
 buffer[1754] = 16'h6147;
 buffer[1755] = 16'h06E1;
 buffer[1756] = 16'h6B8D;
 buffer[1757] = 16'h6103;
 buffer[1758] = 16'h6081;
 buffer[1759] = 16'h6147;
 buffer[1760] = 16'h6A00;
 buffer[1761] = 16'h6181;
 buffer[1762] = 16'h428F;
 buffer[1763] = 16'h6B8D;
 buffer[1764] = 16'h6B8D;
 buffer[1765] = 16'h028F;
 buffer[1766] = 16'h6181;
 buffer[1767] = 16'h6B8D;
 buffer[1768] = 16'h028F;
 buffer[1769] = 16'h0D2E;
 buffer[1770] = 16'h7005;
 buffer[1771] = 16'h7261;
 buffer[1772] = 16'h6573;
 buffer[1773] = 16'h6147;
 buffer[1774] = 16'hFE88;
 buffer[1775] = 16'h6C00;
 buffer[1776] = 16'hFE84;
 buffer[1777] = 16'h6C00;
 buffer[1778] = 16'h6203;
 buffer[1779] = 16'hFE86;
 buffer[1780] = 16'h6C00;
 buffer[1781] = 16'hFE84;
 buffer[1782] = 16'h6C00;
 buffer[1783] = 16'h428F;
 buffer[1784] = 16'h6B8D;
 buffer[1785] = 16'h469B;
 buffer[1786] = 16'hFE84;
 buffer[1787] = 16'h0370;
 buffer[1788] = 16'h0DD4;
 buffer[1789] = 16'h2E82;
 buffer[1790] = 16'h0028;
 buffer[1791] = 16'h8029;
 buffer[1792] = 16'h46ED;
 buffer[1793] = 16'h0519;
 buffer[1794] = 16'h0DFA;
 buffer[1795] = 16'h2881;
 buffer[1796] = 16'h8029;
 buffer[1797] = 16'h46ED;
 buffer[1798] = 16'h0273;
 buffer[1799] = 16'h0E06;
 buffer[1800] = 16'h3C83;
 buffer[1801] = 16'h3E5C;
 buffer[1802] = 16'hFE86;
 buffer[1803] = 16'h6C00;
 buffer[1804] = 16'hFE84;
 buffer[1805] = 16'h6023;
 buffer[1806] = 16'h710F;
 buffer[1807] = 16'h0E10;
 buffer[1808] = 16'h5C81;
 buffer[1809] = 16'hFEB6;
 buffer[1810] = 16'h03BC;
 buffer[1811] = 16'h0E20;
 buffer[1812] = 16'h7704;
 buffer[1813] = 16'h726F;
 buffer[1814] = 16'h0064;
 buffer[1815] = 16'h46ED;
 buffer[1816] = 16'h4394;
 buffer[1817] = 16'h434B;
 buffer[1818] = 16'h05CE;
 buffer[1819] = 16'h0E28;
 buffer[1820] = 16'h7405;
 buffer[1821] = 16'h6B6F;
 buffer[1822] = 16'h6E65;
 buffer[1823] = 16'h435C;
 buffer[1824] = 16'h0717;
 buffer[1825] = 16'h0E38;
 buffer[1826] = 16'h6E05;
 buffer[1827] = 16'h6D61;
 buffer[1828] = 16'h3E65;
 buffer[1829] = 16'h438C;
 buffer[1830] = 16'h801F;
 buffer[1831] = 16'h6303;
 buffer[1832] = 16'h6203;
 buffer[1833] = 16'h039B;
 buffer[1834] = 16'h0E44;
 buffer[1835] = 16'h7305;
 buffer[1836] = 16'h6D61;
 buffer[1837] = 16'h3F65;
 buffer[1838] = 16'h6A00;
 buffer[1839] = 16'h6147;
 buffer[1840] = 16'h073E;
 buffer[1841] = 16'h6181;
 buffer[1842] = 16'h6B81;
 buffer[1843] = 16'h6203;
 buffer[1844] = 16'h417E;
 buffer[1845] = 16'h6181;
 buffer[1846] = 16'h6B81;
 buffer[1847] = 16'h6203;
 buffer[1848] = 16'h417E;
 buffer[1849] = 16'h428F;
 buffer[1850] = 16'h4264;
 buffer[1851] = 16'h273E;
 buffer[1852] = 16'h6B8D;
 buffer[1853] = 16'h710F;
 buffer[1854] = 16'h6B81;
 buffer[1855] = 16'h2744;
 buffer[1856] = 16'h6B8D;
 buffer[1857] = 16'h6A00;
 buffer[1858] = 16'h6147;
 buffer[1859] = 16'h0731;
 buffer[1860] = 16'h6B8D;
 buffer[1861] = 16'h6103;
 buffer[1862] = 16'h8000;
 buffer[1863] = 16'h700C;
 buffer[1864] = 16'h0E56;
 buffer[1865] = 16'h6604;
 buffer[1866] = 16'h6E69;
 buffer[1867] = 16'h0064;
 buffer[1868] = 16'h6180;
 buffer[1869] = 16'h6081;
 buffer[1870] = 16'h417E;
 buffer[1871] = 16'hFE82;
 buffer[1872] = 16'h6023;
 buffer[1873] = 16'h6103;
 buffer[1874] = 16'h6081;
 buffer[1875] = 16'h6C00;
 buffer[1876] = 16'h6147;
 buffer[1877] = 16'h434B;
 buffer[1878] = 16'h6180;
 buffer[1879] = 16'h6C00;
 buffer[1880] = 16'h6081;
 buffer[1881] = 16'h276A;
 buffer[1882] = 16'h6081;
 buffer[1883] = 16'h6C00;
 buffer[1884] = 16'hFF1F;
 buffer[1885] = 16'h6303;
 buffer[1886] = 16'h6B81;
 buffer[1887] = 16'h6503;
 buffer[1888] = 16'h2765;
 buffer[1889] = 16'h434B;
 buffer[1890] = 16'h8000;
 buffer[1891] = 16'h6600;
 buffer[1892] = 16'h0769;
 buffer[1893] = 16'h434B;
 buffer[1894] = 16'hFE82;
 buffer[1895] = 16'h6C00;
 buffer[1896] = 16'h472E;
 buffer[1897] = 16'h076F;
 buffer[1898] = 16'h6B8D;
 buffer[1899] = 16'h6103;
 buffer[1900] = 16'h6180;
 buffer[1901] = 16'h4351;
 buffer[1902] = 16'h718C;
 buffer[1903] = 16'h2774;
 buffer[1904] = 16'h8002;
 buffer[1905] = 16'h4357;
 buffer[1906] = 16'h428F;
 buffer[1907] = 16'h0757;
 buffer[1908] = 16'h6B8D;
 buffer[1909] = 16'h6103;
 buffer[1910] = 16'h6003;
 buffer[1911] = 16'h4351;
 buffer[1912] = 16'h6081;
 buffer[1913] = 16'h4725;
 buffer[1914] = 16'h718C;
 buffer[1915] = 16'h0E92;
 buffer[1916] = 16'h3C07;
 buffer[1917] = 16'h616E;
 buffer[1918] = 16'h656D;
 buffer[1919] = 16'h3E3F;
 buffer[1920] = 16'hFE90;
 buffer[1921] = 16'h6081;
 buffer[1922] = 16'h4383;
 buffer[1923] = 16'h6503;
 buffer[1924] = 16'h2786;
 buffer[1925] = 16'h4351;
 buffer[1926] = 16'h6147;
 buffer[1927] = 16'h6B8D;
 buffer[1928] = 16'h434B;
 buffer[1929] = 16'h6081;
 buffer[1930] = 16'h6147;
 buffer[1931] = 16'h6C00;
 buffer[1932] = 16'h4264;
 buffer[1933] = 16'h2793;
 buffer[1934] = 16'h474C;
 buffer[1935] = 16'h4264;
 buffer[1936] = 16'h2787;
 buffer[1937] = 16'h6B8D;
 buffer[1938] = 16'h710F;
 buffer[1939] = 16'h6B8D;
 buffer[1940] = 16'h6103;
 buffer[1941] = 16'h8000;
 buffer[1942] = 16'h700C;
 buffer[1943] = 16'h0EF8;
 buffer[1944] = 16'h6E05;
 buffer[1945] = 16'h6D61;
 buffer[1946] = 16'h3F65;
 buffer[1947] = 16'hFEB8;
 buffer[1948] = 16'h03BC;
 buffer[1949] = 16'h0F30;
 buffer[1950] = 16'h5E02;
 buffer[1951] = 16'h0068;
 buffer[1952] = 16'h6147;
 buffer[1953] = 16'h6181;
 buffer[1954] = 16'h6B81;
 buffer[1955] = 16'h6803;
 buffer[1956] = 16'h6081;
 buffer[1957] = 16'h27AB;
 buffer[1958] = 16'h8008;
 buffer[1959] = 16'h6081;
 buffer[1960] = 16'h44C7;
 buffer[1961] = 16'h4501;
 buffer[1962] = 16'h44C7;
 buffer[1963] = 16'h6B8D;
 buffer[1964] = 16'h720F;
 buffer[1965] = 16'h0F3C;
 buffer[1966] = 16'h7403;
 buffer[1967] = 16'h7061;
 buffer[1968] = 16'h6081;
 buffer[1969] = 16'h44C7;
 buffer[1970] = 16'h6181;
 buffer[1971] = 16'h418D;
 buffer[1972] = 16'h731C;
 buffer[1973] = 16'h0F5C;
 buffer[1974] = 16'h6B04;
 buffer[1975] = 16'h6174;
 buffer[1976] = 16'h0070;
 buffer[1977] = 16'h6081;
 buffer[1978] = 16'h800D;
 buffer[1979] = 16'h6503;
 buffer[1980] = 16'h27C3;
 buffer[1981] = 16'h8008;
 buffer[1982] = 16'h6503;
 buffer[1983] = 16'h27C2;
 buffer[1984] = 16'h435C;
 buffer[1985] = 16'h07B0;
 buffer[1986] = 16'h07A0;
 buffer[1987] = 16'h6103;
 buffer[1988] = 16'h6003;
 buffer[1989] = 16'h708D;
 buffer[1990] = 16'h0F6C;
 buffer[1991] = 16'h6106;
 buffer[1992] = 16'h6363;
 buffer[1993] = 16'h7065;
 buffer[1994] = 16'h0074;
 buffer[1995] = 16'h6181;
 buffer[1996] = 16'h6203;
 buffer[1997] = 16'h6181;
 buffer[1998] = 16'h4279;
 buffer[1999] = 16'h6503;
 buffer[2000] = 16'h27DC;
 buffer[2001] = 16'h44CC;
 buffer[2002] = 16'h6081;
 buffer[2003] = 16'h435C;
 buffer[2004] = 16'h428F;
 buffer[2005] = 16'h807F;
 buffer[2006] = 16'h6F03;
 buffer[2007] = 16'h27DA;
 buffer[2008] = 16'h47B0;
 buffer[2009] = 16'h07DB;
 buffer[2010] = 16'h47B9;
 buffer[2011] = 16'h07CE;
 buffer[2012] = 16'h6103;
 buffer[2013] = 16'h6181;
 buffer[2014] = 16'h028F;
 buffer[2015] = 16'h0F8E;
 buffer[2016] = 16'h7105;
 buffer[2017] = 16'h6575;
 buffer[2018] = 16'h7972;
 buffer[2019] = 16'hFE88;
 buffer[2020] = 16'h6C00;
 buffer[2021] = 16'h8050;
 buffer[2022] = 16'h47CB;
 buffer[2023] = 16'hFE86;
 buffer[2024] = 16'h6023;
 buffer[2025] = 16'h6103;
 buffer[2026] = 16'h6103;
 buffer[2027] = 16'h8000;
 buffer[2028] = 16'hFE84;
 buffer[2029] = 16'h6023;
 buffer[2030] = 16'h710F;
 buffer[2031] = 16'h0FC0;
 buffer[2032] = 16'h6106;
 buffer[2033] = 16'h6F62;
 buffer[2034] = 16'h7472;
 buffer[2035] = 16'h0032;
 buffer[2036] = 16'h4530;
 buffer[2037] = 16'h710F;
 buffer[2038] = 16'h0FE0;
 buffer[2039] = 16'h6106;
 buffer[2040] = 16'h6F62;
 buffer[2041] = 16'h7472;
 buffer[2042] = 16'h0031;
 buffer[2043] = 16'h4501;
 buffer[2044] = 16'h4542;
 buffer[2045] = 16'h803F;
 buffer[2046] = 16'h44C7;
 buffer[2047] = 16'h4529;
 buffer[2048] = 16'hFE8C;
 buffer[2049] = 16'h43BC;
 buffer[2050] = 16'h07F4;
 buffer[2051] = 16'h0FEE;
 buffer[2052] = 16'h3C49;
 buffer[2053] = 16'h613F;
 buffer[2054] = 16'h6F62;
 buffer[2055] = 16'h7472;
 buffer[2056] = 16'h3E22;
 buffer[2057] = 16'h280C;
 buffer[2058] = 16'h4530;
 buffer[2059] = 16'h07FB;
 buffer[2060] = 16'h07F4;
 buffer[2061] = 16'h1008;
 buffer[2062] = 16'h6606;
 buffer[2063] = 16'h726F;
 buffer[2064] = 16'h6567;
 buffer[2065] = 16'h0074;
 buffer[2066] = 16'h471F;
 buffer[2067] = 16'h479B;
 buffer[2068] = 16'h4264;
 buffer[2069] = 16'h2824;
 buffer[2070] = 16'h4351;
 buffer[2071] = 16'h6081;
 buffer[2072] = 16'hFEAC;
 buffer[2073] = 16'h6023;
 buffer[2074] = 16'h6103;
 buffer[2075] = 16'h6C00;
 buffer[2076] = 16'h6081;
 buffer[2077] = 16'hFE90;
 buffer[2078] = 16'h6023;
 buffer[2079] = 16'h6103;
 buffer[2080] = 16'hFEAE;
 buffer[2081] = 16'h6023;
 buffer[2082] = 16'h6103;
 buffer[2083] = 16'h710F;
 buffer[2084] = 16'h07FB;
 buffer[2085] = 16'h101C;
 buffer[2086] = 16'h240A;
 buffer[2087] = 16'h6E69;
 buffer[2088] = 16'h6574;
 buffer[2089] = 16'h7072;
 buffer[2090] = 16'h6572;
 buffer[2091] = 16'h0074;
 buffer[2092] = 16'h479B;
 buffer[2093] = 16'h4264;
 buffer[2094] = 16'h283C;
 buffer[2095] = 16'h6C00;
 buffer[2096] = 16'h8040;
 buffer[2097] = 16'h6303;
 buffer[2098] = 16'h4809;
 buffer[2099] = 16'h630C;
 buffer[2100] = 16'h6D6F;
 buffer[2101] = 16'h6970;
 buffer[2102] = 16'h656C;
 buffer[2103] = 16'h6F2D;
 buffer[2104] = 16'h6C6E;
 buffer[2105] = 16'h0079;
 buffer[2106] = 16'h0172;
 buffer[2107] = 16'h0840;
 buffer[2108] = 16'h445F;
 buffer[2109] = 16'h283F;
 buffer[2110] = 16'h700C;
 buffer[2111] = 16'h07FB;
 buffer[2112] = 16'h104C;
 buffer[2113] = 16'h5B81;
 buffer[2114] = 16'h9058;
 buffer[2115] = 16'hFE8A;
 buffer[2116] = 16'h6023;
 buffer[2117] = 16'h710F;
 buffer[2118] = 16'h1082;
 buffer[2119] = 16'h2E03;
 buffer[2120] = 16'h6B6F;
 buffer[2121] = 16'h9058;
 buffer[2122] = 16'hFE8A;
 buffer[2123] = 16'h6C00;
 buffer[2124] = 16'h6703;
 buffer[2125] = 16'h2851;
 buffer[2126] = 16'h4547;
 buffer[2127] = 16'h2003;
 buffer[2128] = 16'h6B6F;
 buffer[2129] = 16'h0529;
 buffer[2130] = 16'h108E;
 buffer[2131] = 16'h6504;
 buffer[2132] = 16'h6176;
 buffer[2133] = 16'h006C;
 buffer[2134] = 16'h471F;
 buffer[2135] = 16'h6081;
 buffer[2136] = 16'h417E;
 buffer[2137] = 16'h285D;
 buffer[2138] = 16'hFE8A;
 buffer[2139] = 16'h43BC;
 buffer[2140] = 16'h0856;
 buffer[2141] = 16'h6103;
 buffer[2142] = 16'h0849;
 buffer[2143] = 16'h10A6;
 buffer[2144] = 16'h2445;
 buffer[2145] = 16'h7665;
 buffer[2146] = 16'h6C61;
 buffer[2147] = 16'hFE84;
 buffer[2148] = 16'h6C00;
 buffer[2149] = 16'h6147;
 buffer[2150] = 16'hFE86;
 buffer[2151] = 16'h6C00;
 buffer[2152] = 16'h6147;
 buffer[2153] = 16'hFE88;
 buffer[2154] = 16'h6C00;
 buffer[2155] = 16'h6147;
 buffer[2156] = 16'hFE84;
 buffer[2157] = 16'h8000;
 buffer[2158] = 16'h6180;
 buffer[2159] = 16'h6023;
 buffer[2160] = 16'h6103;
 buffer[2161] = 16'hFE86;
 buffer[2162] = 16'h6023;
 buffer[2163] = 16'h6103;
 buffer[2164] = 16'hFE88;
 buffer[2165] = 16'h6023;
 buffer[2166] = 16'h6103;
 buffer[2167] = 16'h4856;
 buffer[2168] = 16'h6B8D;
 buffer[2169] = 16'hFE88;
 buffer[2170] = 16'h6023;
 buffer[2171] = 16'h6103;
 buffer[2172] = 16'h6B8D;
 buffer[2173] = 16'hFE86;
 buffer[2174] = 16'h6023;
 buffer[2175] = 16'h6103;
 buffer[2176] = 16'h6B8D;
 buffer[2177] = 16'hFE84;
 buffer[2178] = 16'h6023;
 buffer[2179] = 16'h710F;
 buffer[2180] = 16'h10C0;
 buffer[2181] = 16'h7006;
 buffer[2182] = 16'h6572;
 buffer[2183] = 16'h6573;
 buffer[2184] = 16'h0074;
 buffer[2185] = 16'hFF00;
 buffer[2186] = 16'hFE86;
 buffer[2187] = 16'h434B;
 buffer[2188] = 16'h6023;
 buffer[2189] = 16'h710F;
 buffer[2190] = 16'h110A;
 buffer[2191] = 16'h7104;
 buffer[2192] = 16'h6975;
 buffer[2193] = 16'h0074;
 buffer[2194] = 16'h4842;
 buffer[2195] = 16'h47E3;
 buffer[2196] = 16'h4856;
 buffer[2197] = 16'h0893;
 buffer[2198] = 16'h700C;
 buffer[2199] = 16'h111E;
 buffer[2200] = 16'h6105;
 buffer[2201] = 16'h6F62;
 buffer[2202] = 16'h7472;
 buffer[2203] = 16'h6103;
 buffer[2204] = 16'h4889;
 buffer[2205] = 16'h4849;
 buffer[2206] = 16'h0892;
 buffer[2207] = 16'h1130;
 buffer[2208] = 16'h2701;
 buffer[2209] = 16'h471F;
 buffer[2210] = 16'h479B;
 buffer[2211] = 16'h28A5;
 buffer[2212] = 16'h700C;
 buffer[2213] = 16'h07FB;
 buffer[2214] = 16'h1140;
 buffer[2215] = 16'h6105;
 buffer[2216] = 16'h6C6C;
 buffer[2217] = 16'h746F;
 buffer[2218] = 16'h439B;
 buffer[2219] = 16'hFEAC;
 buffer[2220] = 16'h0370;
 buffer[2221] = 16'h114E;
 buffer[2222] = 16'h2C01;
 buffer[2223] = 16'h4394;
 buffer[2224] = 16'h6081;
 buffer[2225] = 16'h434B;
 buffer[2226] = 16'hFEAC;
 buffer[2227] = 16'h6023;
 buffer[2228] = 16'h6103;
 buffer[2229] = 16'h6023;
 buffer[2230] = 16'h710F;
 buffer[2231] = 16'h115C;
 buffer[2232] = 16'h6345;
 buffer[2233] = 16'h6C61;
 buffer[2234] = 16'h2C6C;
 buffer[2235] = 16'h8001;
 buffer[2236] = 16'h6903;
 buffer[2237] = 16'hC000;
 buffer[2238] = 16'h6403;
 buffer[2239] = 16'h08AF;
 buffer[2240] = 16'h1170;
 buffer[2241] = 16'h3F47;
 buffer[2242] = 16'h7262;
 buffer[2243] = 16'h6E61;
 buffer[2244] = 16'h6863;
 buffer[2245] = 16'h8001;
 buffer[2246] = 16'h6903;
 buffer[2247] = 16'hA000;
 buffer[2248] = 16'h6403;
 buffer[2249] = 16'h08AF;
 buffer[2250] = 16'h1182;
 buffer[2251] = 16'h6246;
 buffer[2252] = 16'h6172;
 buffer[2253] = 16'h636E;
 buffer[2254] = 16'h0068;
 buffer[2255] = 16'h8001;
 buffer[2256] = 16'h6903;
 buffer[2257] = 16'h8000;
 buffer[2258] = 16'h6403;
 buffer[2259] = 16'h08AF;
 buffer[2260] = 16'h1196;
 buffer[2261] = 16'h5B89;
 buffer[2262] = 16'h6F63;
 buffer[2263] = 16'h706D;
 buffer[2264] = 16'h6C69;
 buffer[2265] = 16'h5D65;
 buffer[2266] = 16'h48A1;
 buffer[2267] = 16'h08BB;
 buffer[2268] = 16'h11AA;
 buffer[2269] = 16'h6347;
 buffer[2270] = 16'h6D6F;
 buffer[2271] = 16'h6970;
 buffer[2272] = 16'h656C;
 buffer[2273] = 16'h6B8D;
 buffer[2274] = 16'h6081;
 buffer[2275] = 16'h6C00;
 buffer[2276] = 16'h48AF;
 buffer[2277] = 16'h434B;
 buffer[2278] = 16'h6147;
 buffer[2279] = 16'h700C;
 buffer[2280] = 16'h11BA;
 buffer[2281] = 16'h7287;
 buffer[2282] = 16'h6365;
 buffer[2283] = 16'h7275;
 buffer[2284] = 16'h6573;
 buffer[2285] = 16'hFEAE;
 buffer[2286] = 16'h6C00;
 buffer[2287] = 16'h4725;
 buffer[2288] = 16'h08BB;
 buffer[2289] = 16'h11D2;
 buffer[2290] = 16'h7004;
 buffer[2291] = 16'h6369;
 buffer[2292] = 16'h006B;
 buffer[2293] = 16'h6081;
 buffer[2294] = 16'h6410;
 buffer[2295] = 16'h6410;
 buffer[2296] = 16'h80C0;
 buffer[2297] = 16'h6203;
 buffer[2298] = 16'h6147;
 buffer[2299] = 16'h700C;
 buffer[2300] = 16'h11E4;
 buffer[2301] = 16'h6C87;
 buffer[2302] = 16'h7469;
 buffer[2303] = 16'h7265;
 buffer[2304] = 16'h6C61;
 buffer[2305] = 16'h6081;
 buffer[2306] = 16'hFFFF;
 buffer[2307] = 16'h6600;
 buffer[2308] = 16'h6303;
 buffer[2309] = 16'h290D;
 buffer[2310] = 16'h8000;
 buffer[2311] = 16'h6600;
 buffer[2312] = 16'h6503;
 buffer[2313] = 16'h4901;
 buffer[2314] = 16'h48E1;
 buffer[2315] = 16'h6600;
 buffer[2316] = 16'h0911;
 buffer[2317] = 16'hFFFF;
 buffer[2318] = 16'h6600;
 buffer[2319] = 16'h6403;
 buffer[2320] = 16'h08AF;
 buffer[2321] = 16'h700C;
 buffer[2322] = 16'h11FA;
 buffer[2323] = 16'h5B83;
 buffer[2324] = 16'h5D27;
 buffer[2325] = 16'h48A1;
 buffer[2326] = 16'h0901;
 buffer[2327] = 16'h1226;
 buffer[2328] = 16'h2403;
 buffer[2329] = 16'h222C;
 buffer[2330] = 16'h8022;
 buffer[2331] = 16'h46ED;
 buffer[2332] = 16'h4394;
 buffer[2333] = 16'h45CE;
 buffer[2334] = 16'h438C;
 buffer[2335] = 16'h6203;
 buffer[2336] = 16'h439B;
 buffer[2337] = 16'hFEAC;
 buffer[2338] = 16'h6023;
 buffer[2339] = 16'h710F;
 buffer[2340] = 16'h1230;
 buffer[2341] = 16'h66C3;
 buffer[2342] = 16'h726F;
 buffer[2343] = 16'h48E1;
 buffer[2344] = 16'h4112;
 buffer[2345] = 16'h0394;
 buffer[2346] = 16'h124A;
 buffer[2347] = 16'h62C5;
 buffer[2348] = 16'h6765;
 buffer[2349] = 16'h6E69;
 buffer[2350] = 16'h0394;
 buffer[2351] = 16'h1256;
 buffer[2352] = 16'h2846;
 buffer[2353] = 16'h656E;
 buffer[2354] = 16'h7478;
 buffer[2355] = 16'h0029;
 buffer[2356] = 16'h6B8D;
 buffer[2357] = 16'h6B8D;
 buffer[2358] = 16'h4264;
 buffer[2359] = 16'h293D;
 buffer[2360] = 16'h6A00;
 buffer[2361] = 16'h6147;
 buffer[2362] = 16'h6C00;
 buffer[2363] = 16'h6147;
 buffer[2364] = 16'h700C;
 buffer[2365] = 16'h434B;
 buffer[2366] = 16'h6147;
 buffer[2367] = 16'h700C;
 buffer[2368] = 16'h1260;
 buffer[2369] = 16'h6EC4;
 buffer[2370] = 16'h7865;
 buffer[2371] = 16'h0074;
 buffer[2372] = 16'h48E1;
 buffer[2373] = 16'h4934;
 buffer[2374] = 16'h08AF;
 buffer[2375] = 16'h1282;
 buffer[2376] = 16'h2844;
 buffer[2377] = 16'h6F64;
 buffer[2378] = 16'h0029;
 buffer[2379] = 16'h6B8D;
 buffer[2380] = 16'h6081;
 buffer[2381] = 16'h6147;
 buffer[2382] = 16'h6180;
 buffer[2383] = 16'h426B;
 buffer[2384] = 16'h6147;
 buffer[2385] = 16'h6147;
 buffer[2386] = 16'h434B;
 buffer[2387] = 16'h6147;
 buffer[2388] = 16'h700C;
 buffer[2389] = 16'h1290;
 buffer[2390] = 16'h64C2;
 buffer[2391] = 16'h006F;
 buffer[2392] = 16'h48E1;
 buffer[2393] = 16'h494B;
 buffer[2394] = 16'h8000;
 buffer[2395] = 16'h48AF;
 buffer[2396] = 16'h0394;
 buffer[2397] = 16'h12AC;
 buffer[2398] = 16'h2847;
 buffer[2399] = 16'h656C;
 buffer[2400] = 16'h7661;
 buffer[2401] = 16'h2965;
 buffer[2402] = 16'h6B8D;
 buffer[2403] = 16'h6103;
 buffer[2404] = 16'h6B8D;
 buffer[2405] = 16'h6103;
 buffer[2406] = 16'h6B8D;
 buffer[2407] = 16'h710F;
 buffer[2408] = 16'h12BC;
 buffer[2409] = 16'h6CC5;
 buffer[2410] = 16'h6165;
 buffer[2411] = 16'h6576;
 buffer[2412] = 16'h48E1;
 buffer[2413] = 16'h4962;
 buffer[2414] = 16'h700C;
 buffer[2415] = 16'h12D2;
 buffer[2416] = 16'h2846;
 buffer[2417] = 16'h6F6C;
 buffer[2418] = 16'h706F;
 buffer[2419] = 16'h0029;
 buffer[2420] = 16'h6B8D;
 buffer[2421] = 16'h6B8D;
 buffer[2422] = 16'h6310;
 buffer[2423] = 16'h6B8D;
 buffer[2424] = 16'h4279;
 buffer[2425] = 16'h6213;
 buffer[2426] = 16'h2980;
 buffer[2427] = 16'h6147;
 buffer[2428] = 16'h6147;
 buffer[2429] = 16'h6C00;
 buffer[2430] = 16'h6147;
 buffer[2431] = 16'h700C;
 buffer[2432] = 16'h6147;
 buffer[2433] = 16'h6A00;
 buffer[2434] = 16'h6147;
 buffer[2435] = 16'h434B;
 buffer[2436] = 16'h6147;
 buffer[2437] = 16'h700C;
 buffer[2438] = 16'h12E0;
 buffer[2439] = 16'h2848;
 buffer[2440] = 16'h6E75;
 buffer[2441] = 16'h6F6C;
 buffer[2442] = 16'h706F;
 buffer[2443] = 16'h0029;
 buffer[2444] = 16'h6B8D;
 buffer[2445] = 16'h6B8D;
 buffer[2446] = 16'h6103;
 buffer[2447] = 16'h6B8D;
 buffer[2448] = 16'h6103;
 buffer[2449] = 16'h6B8D;
 buffer[2450] = 16'h6103;
 buffer[2451] = 16'h6147;
 buffer[2452] = 16'h700C;
 buffer[2453] = 16'h130E;
 buffer[2454] = 16'h75C6;
 buffer[2455] = 16'h6C6E;
 buffer[2456] = 16'h6F6F;
 buffer[2457] = 16'h0070;
 buffer[2458] = 16'h48E1;
 buffer[2459] = 16'h498C;
 buffer[2460] = 16'h700C;
 buffer[2461] = 16'h132C;
 buffer[2462] = 16'h2845;
 buffer[2463] = 16'h643F;
 buffer[2464] = 16'h296F;
 buffer[2465] = 16'h4279;
 buffer[2466] = 16'h6213;
 buffer[2467] = 16'h29AE;
 buffer[2468] = 16'h6B8D;
 buffer[2469] = 16'h6081;
 buffer[2470] = 16'h6147;
 buffer[2471] = 16'h6180;
 buffer[2472] = 16'h426B;
 buffer[2473] = 16'h6147;
 buffer[2474] = 16'h6147;
 buffer[2475] = 16'h434B;
 buffer[2476] = 16'h6147;
 buffer[2477] = 16'h700C;
 buffer[2478] = 16'h0273;
 buffer[2479] = 16'h700C;
 buffer[2480] = 16'h133C;
 buffer[2481] = 16'h3FC3;
 buffer[2482] = 16'h6F64;
 buffer[2483] = 16'h48E1;
 buffer[2484] = 16'h49A1;
 buffer[2485] = 16'h8000;
 buffer[2486] = 16'h48AF;
 buffer[2487] = 16'h0394;
 buffer[2488] = 16'h1362;
 buffer[2489] = 16'h6CC4;
 buffer[2490] = 16'h6F6F;
 buffer[2491] = 16'h0070;
 buffer[2492] = 16'h48E1;
 buffer[2493] = 16'h4974;
 buffer[2494] = 16'h6081;
 buffer[2495] = 16'h48AF;
 buffer[2496] = 16'h48E1;
 buffer[2497] = 16'h498C;
 buffer[2498] = 16'h4351;
 buffer[2499] = 16'h4394;
 buffer[2500] = 16'h8001;
 buffer[2501] = 16'h6903;
 buffer[2502] = 16'h6180;
 buffer[2503] = 16'h6023;
 buffer[2504] = 16'h710F;
 buffer[2505] = 16'h1372;
 buffer[2506] = 16'h2847;
 buffer[2507] = 16'h6C2B;
 buffer[2508] = 16'h6F6F;
 buffer[2509] = 16'h2970;
 buffer[2510] = 16'h6B8D;
 buffer[2511] = 16'h6180;
 buffer[2512] = 16'h6B8D;
 buffer[2513] = 16'h6B8D;
 buffer[2514] = 16'h4279;
 buffer[2515] = 16'h428F;
 buffer[2516] = 16'h6147;
 buffer[2517] = 16'h8002;
 buffer[2518] = 16'h48F5;
 buffer[2519] = 16'h6B81;
 buffer[2520] = 16'h6203;
 buffer[2521] = 16'h6B81;
 buffer[2522] = 16'h6503;
 buffer[2523] = 16'h6810;
 buffer[2524] = 16'h6010;
 buffer[2525] = 16'h8003;
 buffer[2526] = 16'h48F5;
 buffer[2527] = 16'h6B8D;
 buffer[2528] = 16'h6503;
 buffer[2529] = 16'h6810;
 buffer[2530] = 16'h6010;
 buffer[2531] = 16'h6403;
 buffer[2532] = 16'h29EB;
 buffer[2533] = 16'h6147;
 buffer[2534] = 16'h6203;
 buffer[2535] = 16'h6147;
 buffer[2536] = 16'h6C00;
 buffer[2537] = 16'h6147;
 buffer[2538] = 16'h700C;
 buffer[2539] = 16'h6147;
 buffer[2540] = 16'h6147;
 buffer[2541] = 16'h6103;
 buffer[2542] = 16'h434B;
 buffer[2543] = 16'h6147;
 buffer[2544] = 16'h700C;
 buffer[2545] = 16'h1394;
 buffer[2546] = 16'h2BC5;
 buffer[2547] = 16'h6F6C;
 buffer[2548] = 16'h706F;
 buffer[2549] = 16'h48E1;
 buffer[2550] = 16'h49CE;
 buffer[2551] = 16'h6081;
 buffer[2552] = 16'h48AF;
 buffer[2553] = 16'h48E1;
 buffer[2554] = 16'h498C;
 buffer[2555] = 16'h4351;
 buffer[2556] = 16'h4394;
 buffer[2557] = 16'h8001;
 buffer[2558] = 16'h6903;
 buffer[2559] = 16'h6180;
 buffer[2560] = 16'h6023;
 buffer[2561] = 16'h710F;
 buffer[2562] = 16'h13E4;
 buffer[2563] = 16'h2843;
 buffer[2564] = 16'h2969;
 buffer[2565] = 16'h6B8D;
 buffer[2566] = 16'h6B8D;
 buffer[2567] = 16'h414F;
 buffer[2568] = 16'h6147;
 buffer[2569] = 16'h6147;
 buffer[2570] = 16'h700C;
 buffer[2571] = 16'h1406;
 buffer[2572] = 16'h69C1;
 buffer[2573] = 16'h48E1;
 buffer[2574] = 16'h4A05;
 buffer[2575] = 16'h700C;
 buffer[2576] = 16'h1418;
 buffer[2577] = 16'h75C5;
 buffer[2578] = 16'h746E;
 buffer[2579] = 16'h6C69;
 buffer[2580] = 16'h08C5;
 buffer[2581] = 16'h1422;
 buffer[2582] = 16'h61C5;
 buffer[2583] = 16'h6167;
 buffer[2584] = 16'h6E69;
 buffer[2585] = 16'h08CF;
 buffer[2586] = 16'h142C;
 buffer[2587] = 16'h69C2;
 buffer[2588] = 16'h0066;
 buffer[2589] = 16'h4394;
 buffer[2590] = 16'h8000;
 buffer[2591] = 16'h08C5;
 buffer[2592] = 16'h1436;
 buffer[2593] = 16'h74C4;
 buffer[2594] = 16'h6568;
 buffer[2595] = 16'h006E;
 buffer[2596] = 16'h4394;
 buffer[2597] = 16'h8001;
 buffer[2598] = 16'h6903;
 buffer[2599] = 16'h6181;
 buffer[2600] = 16'h6C00;
 buffer[2601] = 16'h6403;
 buffer[2602] = 16'h6180;
 buffer[2603] = 16'h6023;
 buffer[2604] = 16'h710F;
 buffer[2605] = 16'h1442;
 buffer[2606] = 16'h72C6;
 buffer[2607] = 16'h7065;
 buffer[2608] = 16'h6165;
 buffer[2609] = 16'h0074;
 buffer[2610] = 16'h48CF;
 buffer[2611] = 16'h0A24;
 buffer[2612] = 16'h145C;
 buffer[2613] = 16'h73C4;
 buffer[2614] = 16'h696B;
 buffer[2615] = 16'h0070;
 buffer[2616] = 16'h4394;
 buffer[2617] = 16'h8000;
 buffer[2618] = 16'h08CF;
 buffer[2619] = 16'h146A;
 buffer[2620] = 16'h61C3;
 buffer[2621] = 16'h7466;
 buffer[2622] = 16'h6103;
 buffer[2623] = 16'h4A38;
 buffer[2624] = 16'h492E;
 buffer[2625] = 16'h718C;
 buffer[2626] = 16'h1478;
 buffer[2627] = 16'h65C4;
 buffer[2628] = 16'h736C;
 buffer[2629] = 16'h0065;
 buffer[2630] = 16'h4A38;
 buffer[2631] = 16'h6180;
 buffer[2632] = 16'h0A24;
 buffer[2633] = 16'h1486;
 buffer[2634] = 16'h77C5;
 buffer[2635] = 16'h6968;
 buffer[2636] = 16'h656C;
 buffer[2637] = 16'h4A1D;
 buffer[2638] = 16'h718C;
 buffer[2639] = 16'h1494;
 buffer[2640] = 16'h2846;
 buffer[2641] = 16'h6163;
 buffer[2642] = 16'h6573;
 buffer[2643] = 16'h0029;
 buffer[2644] = 16'h6B8D;
 buffer[2645] = 16'h6180;
 buffer[2646] = 16'h6147;
 buffer[2647] = 16'h6147;
 buffer[2648] = 16'h700C;
 buffer[2649] = 16'h14A0;
 buffer[2650] = 16'h63C4;
 buffer[2651] = 16'h7361;
 buffer[2652] = 16'h0065;
 buffer[2653] = 16'h48E1;
 buffer[2654] = 16'h4A54;
 buffer[2655] = 16'h8030;
 buffer[2656] = 16'h700C;
 buffer[2657] = 16'h14B4;
 buffer[2658] = 16'h2844;
 buffer[2659] = 16'h666F;
 buffer[2660] = 16'h0029;
 buffer[2661] = 16'h6B8D;
 buffer[2662] = 16'h6B81;
 buffer[2663] = 16'h6180;
 buffer[2664] = 16'h6147;
 buffer[2665] = 16'h770F;
 buffer[2666] = 16'h14C4;
 buffer[2667] = 16'h6FC2;
 buffer[2668] = 16'h0066;
 buffer[2669] = 16'h48E1;
 buffer[2670] = 16'h4A65;
 buffer[2671] = 16'h0A1D;
 buffer[2672] = 16'h14D6;
 buffer[2673] = 16'h65C5;
 buffer[2674] = 16'h646E;
 buffer[2675] = 16'h666F;
 buffer[2676] = 16'h4A46;
 buffer[2677] = 16'h8031;
 buffer[2678] = 16'h700C;
 buffer[2679] = 16'h14E2;
 buffer[2680] = 16'h2809;
 buffer[2681] = 16'h6E65;
 buffer[2682] = 16'h6364;
 buffer[2683] = 16'h7361;
 buffer[2684] = 16'h2965;
 buffer[2685] = 16'h6B8D;
 buffer[2686] = 16'h6B8D;
 buffer[2687] = 16'h6103;
 buffer[2688] = 16'h6147;
 buffer[2689] = 16'h700C;
 buffer[2690] = 16'h14F0;
 buffer[2691] = 16'h65C7;
 buffer[2692] = 16'h646E;
 buffer[2693] = 16'h6163;
 buffer[2694] = 16'h6573;
 buffer[2695] = 16'h6081;
 buffer[2696] = 16'h8031;
 buffer[2697] = 16'h6703;
 buffer[2698] = 16'h2A8E;
 buffer[2699] = 16'h6103;
 buffer[2700] = 16'h4A24;
 buffer[2701] = 16'h0A87;
 buffer[2702] = 16'h8030;
 buffer[2703] = 16'h6213;
 buffer[2704] = 16'h4809;
 buffer[2705] = 16'h6213;
 buffer[2706] = 16'h6461;
 buffer[2707] = 16'h6320;
 buffer[2708] = 16'h7361;
 buffer[2709] = 16'h2065;
 buffer[2710] = 16'h6F63;
 buffer[2711] = 16'h736E;
 buffer[2712] = 16'h7274;
 buffer[2713] = 16'h6375;
 buffer[2714] = 16'h2E74;
 buffer[2715] = 16'h48E1;
 buffer[2716] = 16'h4A7D;
 buffer[2717] = 16'h700C;
 buffer[2718] = 16'h1506;
 buffer[2719] = 16'h24C2;
 buffer[2720] = 16'h0022;
 buffer[2721] = 16'h48E1;
 buffer[2722] = 16'h453D;
 buffer[2723] = 16'h091A;
 buffer[2724] = 16'h153E;
 buffer[2725] = 16'h2EC2;
 buffer[2726] = 16'h0022;
 buffer[2727] = 16'h48E1;
 buffer[2728] = 16'h4547;
 buffer[2729] = 16'h091A;
 buffer[2730] = 16'h154A;
 buffer[2731] = 16'h3E05;
 buffer[2732] = 16'h6F62;
 buffer[2733] = 16'h7964;
 buffer[2734] = 16'h034B;
 buffer[2735] = 16'h1556;
 buffer[2736] = 16'h2844;
 buffer[2737] = 16'h6F74;
 buffer[2738] = 16'h0029;
 buffer[2739] = 16'h6B8D;
 buffer[2740] = 16'h6081;
 buffer[2741] = 16'h434B;
 buffer[2742] = 16'h6147;
 buffer[2743] = 16'h6C00;
 buffer[2744] = 16'h6023;
 buffer[2745] = 16'h710F;
 buffer[2746] = 16'h1560;
 buffer[2747] = 16'h74C2;
 buffer[2748] = 16'h006F;
 buffer[2749] = 16'h48E1;
 buffer[2750] = 16'h4AB3;
 buffer[2751] = 16'h48A1;
 buffer[2752] = 16'h4AAE;
 buffer[2753] = 16'h08AF;
 buffer[2754] = 16'h1576;
 buffer[2755] = 16'h2845;
 buffer[2756] = 16'h742B;
 buffer[2757] = 16'h296F;
 buffer[2758] = 16'h6B8D;
 buffer[2759] = 16'h6081;
 buffer[2760] = 16'h434B;
 buffer[2761] = 16'h6147;
 buffer[2762] = 16'h6C00;
 buffer[2763] = 16'h0370;
 buffer[2764] = 16'h1586;
 buffer[2765] = 16'h2BC3;
 buffer[2766] = 16'h6F74;
 buffer[2767] = 16'h48E1;
 buffer[2768] = 16'h4AC6;
 buffer[2769] = 16'h48A1;
 buffer[2770] = 16'h4AAE;
 buffer[2771] = 16'h08AF;
 buffer[2772] = 16'h159A;
 buffer[2773] = 16'h670B;
 buffer[2774] = 16'h7465;
 buffer[2775] = 16'h632D;
 buffer[2776] = 16'h7275;
 buffer[2777] = 16'h6572;
 buffer[2778] = 16'h746E;
 buffer[2779] = 16'hFEA8;
 buffer[2780] = 16'h7C0C;
 buffer[2781] = 16'h15AA;
 buffer[2782] = 16'h730B;
 buffer[2783] = 16'h7465;
 buffer[2784] = 16'h632D;
 buffer[2785] = 16'h7275;
 buffer[2786] = 16'h6572;
 buffer[2787] = 16'h746E;
 buffer[2788] = 16'hFEA8;
 buffer[2789] = 16'h6023;
 buffer[2790] = 16'h710F;
 buffer[2791] = 16'h15BC;
 buffer[2792] = 16'h640B;
 buffer[2793] = 16'h6665;
 buffer[2794] = 16'h6E69;
 buffer[2795] = 16'h7469;
 buffer[2796] = 16'h6F69;
 buffer[2797] = 16'h736E;
 buffer[2798] = 16'hFE90;
 buffer[2799] = 16'h6C00;
 buffer[2800] = 16'h0AE4;
 buffer[2801] = 16'h15D0;
 buffer[2802] = 16'h3F07;
 buffer[2803] = 16'h6E75;
 buffer[2804] = 16'h7169;
 buffer[2805] = 16'h6575;
 buffer[2806] = 16'h6081;
 buffer[2807] = 16'h4ADB;
 buffer[2808] = 16'h474C;
 buffer[2809] = 16'h2B01;
 buffer[2810] = 16'h4547;
 buffer[2811] = 16'h2007;
 buffer[2812] = 16'h6572;
 buffer[2813] = 16'h6564;
 buffer[2814] = 16'h2066;
 buffer[2815] = 16'h6181;
 buffer[2816] = 16'h4542;
 buffer[2817] = 16'h710F;
 buffer[2818] = 16'h15E4;
 buffer[2819] = 16'h3C05;
 buffer[2820] = 16'h2C24;
 buffer[2821] = 16'h3E6E;
 buffer[2822] = 16'h6081;
 buffer[2823] = 16'h417E;
 buffer[2824] = 16'h2B1B;
 buffer[2825] = 16'h4AF6;
 buffer[2826] = 16'h6081;
 buffer[2827] = 16'h438C;
 buffer[2828] = 16'h6203;
 buffer[2829] = 16'h439B;
 buffer[2830] = 16'hFEAC;
 buffer[2831] = 16'h6023;
 buffer[2832] = 16'h6103;
 buffer[2833] = 16'h6081;
 buffer[2834] = 16'hFEAE;
 buffer[2835] = 16'h6023;
 buffer[2836] = 16'h6103;
 buffer[2837] = 16'h4351;
 buffer[2838] = 16'h4ADB;
 buffer[2839] = 16'h6C00;
 buffer[2840] = 16'h6180;
 buffer[2841] = 16'h6023;
 buffer[2842] = 16'h710F;
 buffer[2843] = 16'h6103;
 buffer[2844] = 16'h453D;
 buffer[2845] = 16'h6E04;
 buffer[2846] = 16'h6D61;
 buffer[2847] = 16'h0065;
 buffer[2848] = 16'h07FB;
 buffer[2849] = 16'h1606;
 buffer[2850] = 16'h2403;
 buffer[2851] = 16'h6E2C;
 buffer[2852] = 16'hFEBA;
 buffer[2853] = 16'h03BC;
 buffer[2854] = 16'h1644;
 buffer[2855] = 16'h2408;
 buffer[2856] = 16'h6F63;
 buffer[2857] = 16'h706D;
 buffer[2858] = 16'h6C69;
 buffer[2859] = 16'h0065;
 buffer[2860] = 16'h479B;
 buffer[2861] = 16'h4264;
 buffer[2862] = 16'h2B36;
 buffer[2863] = 16'h6C00;
 buffer[2864] = 16'h8080;
 buffer[2865] = 16'h6303;
 buffer[2866] = 16'h2B35;
 buffer[2867] = 16'h0172;
 buffer[2868] = 16'h0B36;
 buffer[2869] = 16'h08BB;
 buffer[2870] = 16'h445F;
 buffer[2871] = 16'h2B39;
 buffer[2872] = 16'h0901;
 buffer[2873] = 16'h07FB;
 buffer[2874] = 16'h164E;
 buffer[2875] = 16'h6186;
 buffer[2876] = 16'h6F62;
 buffer[2877] = 16'h7472;
 buffer[2878] = 16'h0022;
 buffer[2879] = 16'h48E1;
 buffer[2880] = 16'h4809;
 buffer[2881] = 16'h091A;
 buffer[2882] = 16'h1676;
 buffer[2883] = 16'h3C07;
 buffer[2884] = 16'h766F;
 buffer[2885] = 16'h7265;
 buffer[2886] = 16'h3E74;
 buffer[2887] = 16'hFEAE;
 buffer[2888] = 16'h6C00;
 buffer[2889] = 16'h4ADB;
 buffer[2890] = 16'h6023;
 buffer[2891] = 16'h710F;
 buffer[2892] = 16'h1686;
 buffer[2893] = 16'h6F05;
 buffer[2894] = 16'h6576;
 buffer[2895] = 16'h7472;
 buffer[2896] = 16'hFEBC;
 buffer[2897] = 16'h03BC;
 buffer[2898] = 16'h169A;
 buffer[2899] = 16'h6504;
 buffer[2900] = 16'h6978;
 buffer[2901] = 16'h0074;
 buffer[2902] = 16'h6B8D;
 buffer[2903] = 16'h710F;
 buffer[2904] = 16'h16A6;
 buffer[2905] = 16'h3CC3;
 buffer[2906] = 16'h3E3B;
 buffer[2907] = 16'h48E1;
 buffer[2908] = 16'h4B56;
 buffer[2909] = 16'h4842;
 buffer[2910] = 16'h4B50;
 buffer[2911] = 16'h8000;
 buffer[2912] = 16'h4394;
 buffer[2913] = 16'h6023;
 buffer[2914] = 16'h710F;
 buffer[2915] = 16'h16B2;
 buffer[2916] = 16'h3BC1;
 buffer[2917] = 16'hFEBE;
 buffer[2918] = 16'h03BC;
 buffer[2919] = 16'h16C8;
 buffer[2920] = 16'h5D01;
 buffer[2921] = 16'h9658;
 buffer[2922] = 16'hFE8A;
 buffer[2923] = 16'h6023;
 buffer[2924] = 16'h710F;
 buffer[2925] = 16'h16D0;
 buffer[2926] = 16'h3A01;
 buffer[2927] = 16'h471F;
 buffer[2928] = 16'h4B24;
 buffer[2929] = 16'h0B69;
 buffer[2930] = 16'h16DC;
 buffer[2931] = 16'h6909;
 buffer[2932] = 16'h6D6D;
 buffer[2933] = 16'h6465;
 buffer[2934] = 16'h6169;
 buffer[2935] = 16'h6574;
 buffer[2936] = 16'h8080;
 buffer[2937] = 16'hFEAE;
 buffer[2938] = 16'h6C00;
 buffer[2939] = 16'h6C00;
 buffer[2940] = 16'h6403;
 buffer[2941] = 16'hFEAE;
 buffer[2942] = 16'h6C00;
 buffer[2943] = 16'h6023;
 buffer[2944] = 16'h710F;
 buffer[2945] = 16'h16E6;
 buffer[2946] = 16'h7504;
 buffer[2947] = 16'h6573;
 buffer[2948] = 16'h0072;
 buffer[2949] = 16'h471F;
 buffer[2950] = 16'h4B24;
 buffer[2951] = 16'h4B50;
 buffer[2952] = 16'h48E1;
 buffer[2953] = 16'h41D2;
 buffer[2954] = 16'h08AF;
 buffer[2955] = 16'h1704;
 buffer[2956] = 16'h3C08;
 buffer[2957] = 16'h7263;
 buffer[2958] = 16'h6165;
 buffer[2959] = 16'h6574;
 buffer[2960] = 16'h003E;
 buffer[2961] = 16'h471F;
 buffer[2962] = 16'h4B24;
 buffer[2963] = 16'h4B50;
 buffer[2964] = 16'h838C;
 buffer[2965] = 16'h08BB;
 buffer[2966] = 16'h1718;
 buffer[2967] = 16'h6306;
 buffer[2968] = 16'h6572;
 buffer[2969] = 16'h7461;
 buffer[2970] = 16'h0065;
 buffer[2971] = 16'hFEC0;
 buffer[2972] = 16'h03BC;
 buffer[2973] = 16'h172E;
 buffer[2974] = 16'h7608;
 buffer[2975] = 16'h7261;
 buffer[2976] = 16'h6169;
 buffer[2977] = 16'h6C62;
 buffer[2978] = 16'h0065;
 buffer[2979] = 16'h4B9B;
 buffer[2980] = 16'h8000;
 buffer[2981] = 16'h08AF;
 buffer[2982] = 16'h173C;
 buffer[2983] = 16'h3209;
 buffer[2984] = 16'h6176;
 buffer[2985] = 16'h6972;
 buffer[2986] = 16'h6261;
 buffer[2987] = 16'h656C;
 buffer[2988] = 16'h4B9B;
 buffer[2989] = 16'h8000;
 buffer[2990] = 16'h48AF;
 buffer[2991] = 16'h8001;
 buffer[2992] = 16'h4357;
 buffer[2993] = 16'h08AA;
 buffer[2994] = 16'h174E;
 buffer[2995] = 16'h2847;
 buffer[2996] = 16'h6F64;
 buffer[2997] = 16'h7365;
 buffer[2998] = 16'h293E;
 buffer[2999] = 16'h6B8D;
 buffer[3000] = 16'h8001;
 buffer[3001] = 16'h6903;
 buffer[3002] = 16'h4394;
 buffer[3003] = 16'h8001;
 buffer[3004] = 16'h6903;
 buffer[3005] = 16'hFEAE;
 buffer[3006] = 16'h6C00;
 buffer[3007] = 16'h4725;
 buffer[3008] = 16'h6081;
 buffer[3009] = 16'h434B;
 buffer[3010] = 16'hFFFF;
 buffer[3011] = 16'h6600;
 buffer[3012] = 16'h6403;
 buffer[3013] = 16'h48AF;
 buffer[3014] = 16'h6023;
 buffer[3015] = 16'h6103;
 buffer[3016] = 16'h08AF;
 buffer[3017] = 16'h1766;
 buffer[3018] = 16'h630C;
 buffer[3019] = 16'h6D6F;
 buffer[3020] = 16'h6970;
 buffer[3021] = 16'h656C;
 buffer[3022] = 16'h6F2D;
 buffer[3023] = 16'h6C6E;
 buffer[3024] = 16'h0079;
 buffer[3025] = 16'h8040;
 buffer[3026] = 16'hFEAE;
 buffer[3027] = 16'h6C00;
 buffer[3028] = 16'h6C00;
 buffer[3029] = 16'h6403;
 buffer[3030] = 16'hFEAE;
 buffer[3031] = 16'h6C00;
 buffer[3032] = 16'h6023;
 buffer[3033] = 16'h710F;
 buffer[3034] = 16'h1794;
 buffer[3035] = 16'h6485;
 buffer[3036] = 16'h656F;
 buffer[3037] = 16'h3E73;
 buffer[3038] = 16'h48E1;
 buffer[3039] = 16'h4BB7;
 buffer[3040] = 16'h700C;
 buffer[3041] = 16'h17B6;
 buffer[3042] = 16'h6304;
 buffer[3043] = 16'h6168;
 buffer[3044] = 16'h0072;
 buffer[3045] = 16'h435C;
 buffer[3046] = 16'h4717;
 buffer[3047] = 16'h6310;
 buffer[3048] = 16'h017E;
 buffer[3049] = 16'h17C4;
 buffer[3050] = 16'h5B86;
 buffer[3051] = 16'h6863;
 buffer[3052] = 16'h7261;
 buffer[3053] = 16'h005D;
 buffer[3054] = 16'h4BE5;
 buffer[3055] = 16'h0901;
 buffer[3056] = 16'h17D4;
 buffer[3057] = 16'h6308;
 buffer[3058] = 16'h6E6F;
 buffer[3059] = 16'h7473;
 buffer[3060] = 16'h6E61;
 buffer[3061] = 16'h0074;
 buffer[3062] = 16'h4B9B;
 buffer[3063] = 16'h48AF;
 buffer[3064] = 16'h4BB7;
 buffer[3065] = 16'h7C0C;
 buffer[3066] = 16'h17E2;
 buffer[3067] = 16'h6405;
 buffer[3068] = 16'h6665;
 buffer[3069] = 16'h7265;
 buffer[3070] = 16'h4B9B;
 buffer[3071] = 16'h8000;
 buffer[3072] = 16'h48AF;
 buffer[3073] = 16'h4BB7;
 buffer[3074] = 16'h6C00;
 buffer[3075] = 16'h4264;
 buffer[3076] = 16'h8000;
 buffer[3077] = 16'h6703;
 buffer[3078] = 16'h4809;
 buffer[3079] = 16'h750D;
 buffer[3080] = 16'h696E;
 buffer[3081] = 16'h696E;
 buffer[3082] = 16'h6974;
 buffer[3083] = 16'h6C61;
 buffer[3084] = 16'h7A69;
 buffer[3085] = 16'h6465;
 buffer[3086] = 16'h0172;
 buffer[3087] = 16'h17F6;
 buffer[3088] = 16'h6982;
 buffer[3089] = 16'h0073;
 buffer[3090] = 16'h48A1;
 buffer[3091] = 16'h4AAE;
 buffer[3092] = 16'h6023;
 buffer[3093] = 16'h710F;
 buffer[3094] = 16'h1820;
 buffer[3095] = 16'h2E03;
 buffer[3096] = 16'h6469;
 buffer[3097] = 16'h4264;
 buffer[3098] = 16'h2C1F;
 buffer[3099] = 16'h438C;
 buffer[3100] = 16'h801F;
 buffer[3101] = 16'h6303;
 buffer[3102] = 16'h0519;
 buffer[3103] = 16'h4529;
 buffer[3104] = 16'h4547;
 buffer[3105] = 16'h7B08;
 buffer[3106] = 16'h6F6E;
 buffer[3107] = 16'h616E;
 buffer[3108] = 16'h656D;
 buffer[3109] = 16'h007D;
 buffer[3110] = 16'h700C;
 buffer[3111] = 16'h182E;
 buffer[3112] = 16'h7708;
 buffer[3113] = 16'h726F;
 buffer[3114] = 16'h6C64;
 buffer[3115] = 16'h7369;
 buffer[3116] = 16'h0074;
 buffer[3117] = 16'h43AA;
 buffer[3118] = 16'h4394;
 buffer[3119] = 16'h8000;
 buffer[3120] = 16'h48AF;
 buffer[3121] = 16'h6081;
 buffer[3122] = 16'hFEA8;
 buffer[3123] = 16'h434B;
 buffer[3124] = 16'h6081;
 buffer[3125] = 16'h6C00;
 buffer[3126] = 16'h48AF;
 buffer[3127] = 16'h6023;
 buffer[3128] = 16'h6103;
 buffer[3129] = 16'h8000;
 buffer[3130] = 16'h08AF;
 buffer[3131] = 16'h1850;
 buffer[3132] = 16'h6F06;
 buffer[3133] = 16'h6472;
 buffer[3134] = 16'h7265;
 buffer[3135] = 16'h0040;
 buffer[3136] = 16'h6081;
 buffer[3137] = 16'h6C00;
 buffer[3138] = 16'h6081;
 buffer[3139] = 16'h2C4A;
 buffer[3140] = 16'h6147;
 buffer[3141] = 16'h434B;
 buffer[3142] = 16'h4C40;
 buffer[3143] = 16'h6B8D;
 buffer[3144] = 16'h6180;
 buffer[3145] = 16'h731C;
 buffer[3146] = 16'h700F;
 buffer[3147] = 16'h1878;
 buffer[3148] = 16'h6709;
 buffer[3149] = 16'h7465;
 buffer[3150] = 16'h6F2D;
 buffer[3151] = 16'h6472;
 buffer[3152] = 16'h7265;
 buffer[3153] = 16'hFE90;
 buffer[3154] = 16'h0C40;
 buffer[3155] = 16'h1898;
 buffer[3156] = 16'h3E04;
 buffer[3157] = 16'h6977;
 buffer[3158] = 16'h0064;
 buffer[3159] = 16'h034B;
 buffer[3160] = 16'h18A8;
 buffer[3161] = 16'h2E04;
 buffer[3162] = 16'h6977;
 buffer[3163] = 16'h0064;
 buffer[3164] = 16'h4501;
 buffer[3165] = 16'h6081;
 buffer[3166] = 16'h4C57;
 buffer[3167] = 16'h434B;
 buffer[3168] = 16'h6C00;
 buffer[3169] = 16'h4264;
 buffer[3170] = 16'h2C65;
 buffer[3171] = 16'h4C19;
 buffer[3172] = 16'h710F;
 buffer[3173] = 16'h8000;
 buffer[3174] = 16'h0556;
 buffer[3175] = 16'h18B2;
 buffer[3176] = 16'h2104;
 buffer[3177] = 16'h6977;
 buffer[3178] = 16'h0064;
 buffer[3179] = 16'h4C57;
 buffer[3180] = 16'h434B;
 buffer[3181] = 16'hFEAE;
 buffer[3182] = 16'h6C00;
 buffer[3183] = 16'h6180;
 buffer[3184] = 16'h6023;
 buffer[3185] = 16'h710F;
 buffer[3186] = 16'h18D0;
 buffer[3187] = 16'h7604;
 buffer[3188] = 16'h636F;
 buffer[3189] = 16'h0073;
 buffer[3190] = 16'h4529;
 buffer[3191] = 16'h4547;
 buffer[3192] = 16'h7605;
 buffer[3193] = 16'h636F;
 buffer[3194] = 16'h3A73;
 buffer[3195] = 16'hFEA8;
 buffer[3196] = 16'h434B;
 buffer[3197] = 16'h6C00;
 buffer[3198] = 16'h4264;
 buffer[3199] = 16'h2C84;
 buffer[3200] = 16'h6081;
 buffer[3201] = 16'h4C5C;
 buffer[3202] = 16'h4C57;
 buffer[3203] = 16'h0C7D;
 buffer[3204] = 16'h700C;
 buffer[3205] = 16'h18E6;
 buffer[3206] = 16'h6F05;
 buffer[3207] = 16'h6472;
 buffer[3208] = 16'h7265;
 buffer[3209] = 16'h4529;
 buffer[3210] = 16'h4547;
 buffer[3211] = 16'h7307;
 buffer[3212] = 16'h6165;
 buffer[3213] = 16'h6372;
 buffer[3214] = 16'h3A68;
 buffer[3215] = 16'h4C51;
 buffer[3216] = 16'h4264;
 buffer[3217] = 16'h2C96;
 buffer[3218] = 16'h6180;
 buffer[3219] = 16'h4C5C;
 buffer[3220] = 16'h6A00;
 buffer[3221] = 16'h0C90;
 buffer[3222] = 16'h4529;
 buffer[3223] = 16'h4547;
 buffer[3224] = 16'h6407;
 buffer[3225] = 16'h6665;
 buffer[3226] = 16'h6E69;
 buffer[3227] = 16'h3A65;
 buffer[3228] = 16'h4ADB;
 buffer[3229] = 16'h0C5C;
 buffer[3230] = 16'h190C;
 buffer[3231] = 16'h7309;
 buffer[3232] = 16'h7465;
 buffer[3233] = 16'h6F2D;
 buffer[3234] = 16'h6472;
 buffer[3235] = 16'h7265;
 buffer[3236] = 16'h6081;
 buffer[3237] = 16'h8000;
 buffer[3238] = 16'h6600;
 buffer[3239] = 16'h6703;
 buffer[3240] = 16'h2CAC;
 buffer[3241] = 16'h6103;
 buffer[3242] = 16'hFEA2;
 buffer[3243] = 16'h8001;
 buffer[3244] = 16'h8008;
 buffer[3245] = 16'h6181;
 buffer[3246] = 16'h6F03;
 buffer[3247] = 16'h4809;
 buffer[3248] = 16'h6F12;
 buffer[3249] = 16'h6576;
 buffer[3250] = 16'h2072;
 buffer[3251] = 16'h6973;
 buffer[3252] = 16'h657A;
 buffer[3253] = 16'h6F20;
 buffer[3254] = 16'h2066;
 buffer[3255] = 16'h7623;
 buffer[3256] = 16'h636F;
 buffer[3257] = 16'h0073;
 buffer[3258] = 16'hFE90;
 buffer[3259] = 16'h6180;
 buffer[3260] = 16'h6081;
 buffer[3261] = 16'h2CC7;
 buffer[3262] = 16'h6147;
 buffer[3263] = 16'h6180;
 buffer[3264] = 16'h6181;
 buffer[3265] = 16'h6023;
 buffer[3266] = 16'h6103;
 buffer[3267] = 16'h434B;
 buffer[3268] = 16'h6B8D;
 buffer[3269] = 16'h6A00;
 buffer[3270] = 16'h0CBC;
 buffer[3271] = 16'h6180;
 buffer[3272] = 16'h6023;
 buffer[3273] = 16'h710F;
 buffer[3274] = 16'h193E;
 buffer[3275] = 16'h6F04;
 buffer[3276] = 16'h6C6E;
 buffer[3277] = 16'h0079;
 buffer[3278] = 16'h8000;
 buffer[3279] = 16'h6600;
 buffer[3280] = 16'h0CA4;
 buffer[3281] = 16'h1996;
 buffer[3282] = 16'h6104;
 buffer[3283] = 16'h736C;
 buffer[3284] = 16'h006F;
 buffer[3285] = 16'h4C51;
 buffer[3286] = 16'h6181;
 buffer[3287] = 16'h6180;
 buffer[3288] = 16'h6310;
 buffer[3289] = 16'h0CA4;
 buffer[3290] = 16'h19A4;
 buffer[3291] = 16'h7008;
 buffer[3292] = 16'h6572;
 buffer[3293] = 16'h6976;
 buffer[3294] = 16'h756F;
 buffer[3295] = 16'h0073;
 buffer[3296] = 16'h4C51;
 buffer[3297] = 16'h6180;
 buffer[3298] = 16'h6103;
 buffer[3299] = 16'h6A00;
 buffer[3300] = 16'h0CA4;
 buffer[3301] = 16'h19B6;
 buffer[3302] = 16'h3E04;
 buffer[3303] = 16'h6F76;
 buffer[3304] = 16'h0063;
 buffer[3305] = 16'h4B9B;
 buffer[3306] = 16'h6081;
 buffer[3307] = 16'h48AF;
 buffer[3308] = 16'h4C6B;
 buffer[3309] = 16'h4BB7;
 buffer[3310] = 16'h6C00;
 buffer[3311] = 16'h6147;
 buffer[3312] = 16'h4C51;
 buffer[3313] = 16'h6180;
 buffer[3314] = 16'h6103;
 buffer[3315] = 16'h6B8D;
 buffer[3316] = 16'h6180;
 buffer[3317] = 16'h0CA4;
 buffer[3318] = 16'h19CC;
 buffer[3319] = 16'h7705;
 buffer[3320] = 16'h6469;
 buffer[3321] = 16'h666F;
 buffer[3322] = 16'h48A1;
 buffer[3323] = 16'h4AAE;
 buffer[3324] = 16'h7C0C;
 buffer[3325] = 16'h19EE;
 buffer[3326] = 16'h760A;
 buffer[3327] = 16'h636F;
 buffer[3328] = 16'h6261;
 buffer[3329] = 16'h6C75;
 buffer[3330] = 16'h7261;
 buffer[3331] = 16'h0079;
 buffer[3332] = 16'h4C2D;
 buffer[3333] = 16'h0CE9;
 buffer[3334] = 16'h19FC;
 buffer[3335] = 16'h5F05;
 buffer[3336] = 16'h7974;
 buffer[3337] = 16'h6570;
 buffer[3338] = 16'h6147;
 buffer[3339] = 16'h0D0F;
 buffer[3340] = 16'h438C;
 buffer[3341] = 16'h4362;
 buffer[3342] = 16'h44C7;
 buffer[3343] = 16'h6B81;
 buffer[3344] = 16'h2D15;
 buffer[3345] = 16'h6B8D;
 buffer[3346] = 16'h6A00;
 buffer[3347] = 16'h6147;
 buffer[3348] = 16'h0D0C;
 buffer[3349] = 16'h6B8D;
 buffer[3350] = 16'h6103;
 buffer[3351] = 16'h710F;
 buffer[3352] = 16'h1A0E;
 buffer[3353] = 16'h6403;
 buffer[3354] = 16'h2B6D;
 buffer[3355] = 16'h6181;
 buffer[3356] = 16'h8004;
 buffer[3357] = 16'h4556;
 buffer[3358] = 16'h4501;
 buffer[3359] = 16'h6147;
 buffer[3360] = 16'h0D24;
 buffer[3361] = 16'h438C;
 buffer[3362] = 16'h8003;
 buffer[3363] = 16'h4556;
 buffer[3364] = 16'h6B81;
 buffer[3365] = 16'h2D2A;
 buffer[3366] = 16'h6B8D;
 buffer[3367] = 16'h6A00;
 buffer[3368] = 16'h6147;
 buffer[3369] = 16'h0D21;
 buffer[3370] = 16'h6B8D;
 buffer[3371] = 16'h710F;
 buffer[3372] = 16'h1A32;
 buffer[3373] = 16'h6404;
 buffer[3374] = 16'h6D75;
 buffer[3375] = 16'h0070;
 buffer[3376] = 16'hFE80;
 buffer[3377] = 16'h6C00;
 buffer[3378] = 16'h6147;
 buffer[3379] = 16'h4432;
 buffer[3380] = 16'h8010;
 buffer[3381] = 16'h4305;
 buffer[3382] = 16'h6147;
 buffer[3383] = 16'h4529;
 buffer[3384] = 16'h8010;
 buffer[3385] = 16'h4279;
 buffer[3386] = 16'h4D1B;
 buffer[3387] = 16'h4155;
 buffer[3388] = 16'h8002;
 buffer[3389] = 16'h4508;
 buffer[3390] = 16'h4D0A;
 buffer[3391] = 16'h6B81;
 buffer[3392] = 16'h2D45;
 buffer[3393] = 16'h6B8D;
 buffer[3394] = 16'h6A00;
 buffer[3395] = 16'h6147;
 buffer[3396] = 16'h0D37;
 buffer[3397] = 16'h6B8D;
 buffer[3398] = 16'h6103;
 buffer[3399] = 16'h6103;
 buffer[3400] = 16'h6B8D;
 buffer[3401] = 16'hFE80;
 buffer[3402] = 16'h6023;
 buffer[3403] = 16'h710F;
 buffer[3404] = 16'h1A5A;
 buffer[3405] = 16'h2E02;
 buffer[3406] = 16'h0073;
 buffer[3407] = 16'h4529;
 buffer[3408] = 16'h416A;
 buffer[3409] = 16'h6A00;
 buffer[3410] = 16'h800F;
 buffer[3411] = 16'h6303;
 buffer[3412] = 16'h6147;
 buffer[3413] = 16'h6B81;
 buffer[3414] = 16'h48F5;
 buffer[3415] = 16'h4569;
 buffer[3416] = 16'h6B81;
 buffer[3417] = 16'h2D5E;
 buffer[3418] = 16'h6B8D;
 buffer[3419] = 16'h6A00;
 buffer[3420] = 16'h6147;
 buffer[3421] = 16'h0D55;
 buffer[3422] = 16'h6B8D;
 buffer[3423] = 16'h6103;
 buffer[3424] = 16'h4547;
 buffer[3425] = 16'h3C04;
 buffer[3426] = 16'h6F74;
 buffer[3427] = 16'h0073;
 buffer[3428] = 16'h700C;
 buffer[3429] = 16'h1A9A;
 buffer[3430] = 16'h2807;
 buffer[3431] = 16'h6E3E;
 buffer[3432] = 16'h6D61;
 buffer[3433] = 16'h2965;
 buffer[3434] = 16'h6C00;
 buffer[3435] = 16'h4264;
 buffer[3436] = 16'h2D74;
 buffer[3437] = 16'h4279;
 buffer[3438] = 16'h4725;
 buffer[3439] = 16'h6503;
 buffer[3440] = 16'h2D73;
 buffer[3441] = 16'h4351;
 buffer[3442] = 16'h0D6A;
 buffer[3443] = 16'h700F;
 buffer[3444] = 16'h6103;
 buffer[3445] = 16'h8000;
 buffer[3446] = 16'h700C;
 buffer[3447] = 16'h1ACC;
 buffer[3448] = 16'h3E05;
 buffer[3449] = 16'h616E;
 buffer[3450] = 16'h656D;
 buffer[3451] = 16'h6147;
 buffer[3452] = 16'h4C51;
 buffer[3453] = 16'h4264;
 buffer[3454] = 16'h2D97;
 buffer[3455] = 16'h6180;
 buffer[3456] = 16'h6B81;
 buffer[3457] = 16'h6180;
 buffer[3458] = 16'h4D6A;
 buffer[3459] = 16'h4264;
 buffer[3460] = 16'h2D95;
 buffer[3461] = 16'h6147;
 buffer[3462] = 16'h6A00;
 buffer[3463] = 16'h6147;
 buffer[3464] = 16'h0D8A;
 buffer[3465] = 16'h6103;
 buffer[3466] = 16'h6B81;
 buffer[3467] = 16'h2D90;
 buffer[3468] = 16'h6B8D;
 buffer[3469] = 16'h6A00;
 buffer[3470] = 16'h6147;
 buffer[3471] = 16'h0D89;
 buffer[3472] = 16'h6B8D;
 buffer[3473] = 16'h6103;
 buffer[3474] = 16'h6B8D;
 buffer[3475] = 16'h6B8D;
 buffer[3476] = 16'h710F;
 buffer[3477] = 16'h6A00;
 buffer[3478] = 16'h0D7D;
 buffer[3479] = 16'h6B8D;
 buffer[3480] = 16'h6103;
 buffer[3481] = 16'h8000;
 buffer[3482] = 16'h700C;
 buffer[3483] = 16'h1AF0;
 buffer[3484] = 16'h7303;
 buffer[3485] = 16'h6565;
 buffer[3486] = 16'h48A1;
 buffer[3487] = 16'h4529;
 buffer[3488] = 16'h6081;
 buffer[3489] = 16'h6C00;
 buffer[3490] = 16'h4264;
 buffer[3491] = 16'hF00C;
 buffer[3492] = 16'h6503;
 buffer[3493] = 16'h2DB7;
 buffer[3494] = 16'hBFFF;
 buffer[3495] = 16'h6303;
 buffer[3496] = 16'h8001;
 buffer[3497] = 16'h6D03;
 buffer[3498] = 16'h4D7B;
 buffer[3499] = 16'h4264;
 buffer[3500] = 16'h2DB0;
 buffer[3501] = 16'h4501;
 buffer[3502] = 16'h4C19;
 buffer[3503] = 16'h0DB5;
 buffer[3504] = 16'h6081;
 buffer[3505] = 16'h6C00;
 buffer[3506] = 16'hFFFF;
 buffer[3507] = 16'h6303;
 buffer[3508] = 16'h4562;
 buffer[3509] = 16'h434B;
 buffer[3510] = 16'h0DA0;
 buffer[3511] = 16'h0273;
 buffer[3512] = 16'h1B38;
 buffer[3513] = 16'h2807;
 buffer[3514] = 16'h6F77;
 buffer[3515] = 16'h6472;
 buffer[3516] = 16'h2973;
 buffer[3517] = 16'h4529;
 buffer[3518] = 16'h6C00;
 buffer[3519] = 16'h4264;
 buffer[3520] = 16'h2DC6;
 buffer[3521] = 16'h6081;
 buffer[3522] = 16'h4C19;
 buffer[3523] = 16'h4501;
 buffer[3524] = 16'h4351;
 buffer[3525] = 16'h0DBE;
 buffer[3526] = 16'h700C;
 buffer[3527] = 16'h1B72;
 buffer[3528] = 16'h7705;
 buffer[3529] = 16'h726F;
 buffer[3530] = 16'h7364;
 buffer[3531] = 16'h4C51;
 buffer[3532] = 16'h4264;
 buffer[3533] = 16'h2DD9;
 buffer[3534] = 16'h6180;
 buffer[3535] = 16'h4529;
 buffer[3536] = 16'h4529;
 buffer[3537] = 16'h4547;
 buffer[3538] = 16'h3A01;
 buffer[3539] = 16'h6081;
 buffer[3540] = 16'h4C5C;
 buffer[3541] = 16'h4529;
 buffer[3542] = 16'h4DBD;
 buffer[3543] = 16'h6A00;
 buffer[3544] = 16'h0DCC;
 buffer[3545] = 16'h700C;
 buffer[3546] = 16'h1B90;
 buffer[3547] = 16'h7603;
 buffer[3548] = 16'h7265;
 buffer[3549] = 16'h8001;
 buffer[3550] = 16'h8100;
 buffer[3551] = 16'h4329;
 buffer[3552] = 16'h8005;
 buffer[3553] = 16'h720F;
 buffer[3554] = 16'h1BB6;
 buffer[3555] = 16'h6802;
 buffer[3556] = 16'h0069;
 buffer[3557] = 16'h4529;
 buffer[3558] = 16'h4547;
 buffer[3559] = 16'h650C;
 buffer[3560] = 16'h6F66;
 buffer[3561] = 16'h7472;
 buffer[3562] = 16'h2068;
 buffer[3563] = 16'h316A;
 buffer[3564] = 16'h202B;
 buffer[3565] = 16'h0076;
 buffer[3566] = 16'hFE80;
 buffer[3567] = 16'h6C00;
 buffer[3568] = 16'h4432;
 buffer[3569] = 16'h4DDD;
 buffer[3570] = 16'h43F4;
 buffer[3571] = 16'h4406;
 buffer[3572] = 16'h4406;
 buffer[3573] = 16'h802E;
 buffer[3574] = 16'h43FC;
 buffer[3575] = 16'h4406;
 buffer[3576] = 16'h441E;
 buffer[3577] = 16'h4519;
 buffer[3578] = 16'hFE80;
 buffer[3579] = 16'h6023;
 buffer[3580] = 16'h6103;
 buffer[3581] = 16'h0529;
 buffer[3582] = 16'h1BC6;
 buffer[3583] = 16'h6304;
 buffer[3584] = 16'h6C6F;
 buffer[3585] = 16'h0064;
 buffer[3586] = 16'h8002;
 buffer[3587] = 16'hFE80;
 buffer[3588] = 16'h8042;
 buffer[3589] = 16'h45B7;
 buffer[3590] = 16'h4889;
 buffer[3591] = 16'hFEA2;
 buffer[3592] = 16'h6081;
 buffer[3593] = 16'hFE90;
 buffer[3594] = 16'h6023;
 buffer[3595] = 16'h6103;
 buffer[3596] = 16'h6081;
 buffer[3597] = 16'hFEA8;
 buffer[3598] = 16'h4379;
 buffer[3599] = 16'h4B50;
 buffer[3600] = 16'hC000;
 buffer[3601] = 16'h434B;
 buffer[3602] = 16'h6081;
 buffer[3603] = 16'h4351;
 buffer[3604] = 16'h6C00;
 buffer[3605] = 16'h4863;
 buffer[3606] = 16'hFEB4;
 buffer[3607] = 16'h43BC;
 buffer[3608] = 16'h4892;
 buffer[3609] = 16'h0E02;
end

endmodule

module M_main_mem_ram(
input      [0:0]             in_ram_wenable0,
input       [15:0]     in_ram_wdata0,
input      [14:0]                in_ram_addr0,
input      [0:0]             in_ram_wenable1,
input      [15:0]                 in_ram_wdata1,
input      [14:0]                in_ram_addr1,
output reg  [15:0]     out_ram_rdata0,
output reg  [15:0]     out_ram_rdata1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[32767:0];
always @(posedge clock0) begin
  if (in_ram_wenable0) begin
    buffer[in_ram_addr0] <= in_ram_wdata0;
  end else begin
    out_ram_rdata0 <= buffer[in_ram_addr0];
  end
end
always @(posedge clock1) begin
  if (in_ram_wenable1) begin
    buffer[in_ram_addr1] <= in_ram_wdata1;
  end else begin
    out_ram_rdata1 <= buffer[in_ram_addr1];
  end
end

endmodule

module M_main_mem_uartInBuffer(
input      [0:0]             in_uartInBuffer_wenable0,
input       [7:0]     in_uartInBuffer_wdata0,
input      [8:0]                in_uartInBuffer_addr0,
input      [0:0]             in_uartInBuffer_wenable1,
input      [7:0]                 in_uartInBuffer_wdata1,
input      [8:0]                in_uartInBuffer_addr1,
output reg  [7:0]     out_uartInBuffer_rdata0,
output reg  [7:0]     out_uartInBuffer_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[511:0];
always @(posedge clock0) begin
  if (in_uartInBuffer_wenable0) begin
    buffer[in_uartInBuffer_addr0] <= in_uartInBuffer_wdata0;
  end else begin
    out_uartInBuffer_rdata0 <= buffer[in_uartInBuffer_addr0];
  end
end
always @(posedge clock1) begin
  if (in_uartInBuffer_wenable1) begin
    buffer[in_uartInBuffer_addr1] <= in_uartInBuffer_wdata1;
  end else begin
    out_uartInBuffer_rdata1 <= buffer[in_uartInBuffer_addr1];
  end
end

endmodule

module M_main_mem_uartOutBuffer(
input      [0:0]             in_uartOutBuffer_wenable0,
input       [7:0]     in_uartOutBuffer_wdata0,
input      [8:0]                in_uartOutBuffer_addr0,
input      [0:0]             in_uartOutBuffer_wenable1,
input      [7:0]                 in_uartOutBuffer_wdata1,
input      [8:0]                in_uartOutBuffer_addr1,
output reg  [7:0]     out_uartOutBuffer_rdata0,
output reg  [7:0]     out_uartOutBuffer_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[511:0];
always @(posedge clock0) begin
  if (in_uartOutBuffer_wenable0) begin
    buffer[in_uartOutBuffer_addr0] <= in_uartOutBuffer_wdata0;
  end else begin
    out_uartOutBuffer_rdata0 <= buffer[in_uartOutBuffer_addr0];
  end
end
always @(posedge clock1) begin
  if (in_uartOutBuffer_wenable1) begin
    buffer[in_uartOutBuffer_addr1] <= in_uartOutBuffer_wdata1;
  end else begin
    out_uartOutBuffer_rdata1 <= buffer[in_uartOutBuffer_addr1];
  end
end

endmodule

module M_main (
in_buttons,
in_uart_tx_busy,
in_uart_rx_data,
in_uart_rx_valid,
in_timer1hz,
out_led,
out_uart_tx_data,
out_uart_tx_valid,
in_run,
out_done,
reset,
clock
);
input  [3:0] in_buttons;
input  [0:0] in_uart_tx_busy;
input  [7:0] in_uart_rx_data;
input  [0:0] in_uart_rx_valid;
input  [15:0] in_timer1hz;
output  [7:0] out_led;
output  [7:0] out_uart_tx_data;
output  [0:0] out_uart_tx_valid;
input in_run;
output out_done;
input reset;
input clock;
wire  [15:0] _w_mem_dstack_rdata;
wire  [15:0] _w_mem_rstack_rdata;
wire  [15:0] _w_mem_rom_rdata;
wire  [15:0] _w_mem_ram_rdata0;
wire  [15:0] _w_mem_ram_rdata1;
wire  [7:0] _w_mem_uartInBuffer_rdata0;
wire  [7:0] _w_mem_uartInBuffer_rdata1;
wire  [7:0] _w_mem_uartOutBuffer_rdata0;
wire  [7:0] _w_mem_uartOutBuffer_rdata1;
wire  [15:0] _c_ram_wdata1;
assign _c_ram_wdata1 = 0;
wire  [7:0] _c_uartInBuffer_wdata0;
assign _c_uartInBuffer_wdata0 = 0;
wire  [7:0] _c_uartOutBuffer_wdata0;
assign _c_uartOutBuffer_wdata0 = 0;
wire  [15:0] _w_immediate;
wire  [0:0] _w_is_alu;
wire  [0:0] _w_is_call;
wire  [0:0] _w_is_lit;
wire  [0:0] _w_dstackWrite;
wire  [0:0] _w_rstackWrite;
wire  [7:0] _w_ddelta;
wire  [7:0] _w_rdelta;
wire  [12:0] _w_pcPlusOne;

reg  [15:0] _d_instruction;
reg  [15:0] _q_instruction;
reg  [12:0] _d_pc;
reg  [12:0] _q_pc;
reg  [12:0] _d_newPC;
reg  [12:0] _q_newPC;
reg  [0:0] _d_dstack_wenable;
reg  [0:0] _q_dstack_wenable;
reg  [15:0] _d_dstack_wdata;
reg  [15:0] _q_dstack_wdata;
reg  [7:0] _d_dstack_addr;
reg  [7:0] _q_dstack_addr;
reg  [15:0] _d_stackTop;
reg  [15:0] _q_stackTop;
reg  [7:0] _d_dsp;
reg  [7:0] _q_dsp;
reg  [7:0] _d_newDSP;
reg  [7:0] _q_newDSP;
reg  [15:0] _d_newStackTop;
reg  [15:0] _q_newStackTop;
reg  [0:0] _d_rstack_wenable;
reg  [0:0] _q_rstack_wenable;
reg  [15:0] _d_rstack_wdata;
reg  [15:0] _q_rstack_wdata;
reg  [7:0] _d_rstack_addr;
reg  [7:0] _q_rstack_addr;
reg  [7:0] _d_rsp;
reg  [7:0] _q_rsp;
reg  [7:0] _d_newRSP;
reg  [7:0] _q_newRSP;
reg  [15:0] _d_rstackWData;
reg  [15:0] _q_rstackWData;
reg  [15:0] _d_stackNext;
reg  [15:0] _q_stackNext;
reg  [15:0] _d_rStackTop;
reg  [15:0] _q_rStackTop;
reg  [15:0] _d_memoryInput;
reg  [15:0] _q_memoryInput;
reg  [11:0] _d_rom_addr;
reg  [11:0] _q_rom_addr;
reg  [0:0] _d_ram_wenable0;
reg  [0:0] _q_ram_wenable0;
reg  [15:0] _d_ram_wdata0;
reg  [15:0] _q_ram_wdata0;
reg  [14:0] _d_ram_addr0;
reg  [14:0] _q_ram_addr0;
reg  [0:0] _d_ram_wenable1;
reg  [0:0] _q_ram_wenable1;
reg  [14:0] _d_ram_addr1;
reg  [14:0] _q_ram_addr1;
reg  [19:0] _d_CYCLE;
reg  [19:0] _q_CYCLE;
reg  [1:0] _d_INIT;
reg  [1:0] _q_INIT;
reg  [15:0] _d_copyaddress;
reg  [15:0] _q_copyaddress;
reg  [15:0] _d_bramREAD;
reg  [15:0] _q_bramREAD;
reg  [0:0] _d_uartInBuffer_wenable0;
reg  [0:0] _q_uartInBuffer_wenable0;
reg  [8:0] _d_uartInBuffer_addr0;
reg  [8:0] _q_uartInBuffer_addr0;
reg  [0:0] _d_uartInBuffer_wenable1;
reg  [0:0] _q_uartInBuffer_wenable1;
reg  [7:0] _d_uartInBuffer_wdata1;
reg  [7:0] _q_uartInBuffer_wdata1;
reg  [8:0] _d_uartInBuffer_addr1;
reg  [8:0] _q_uartInBuffer_addr1;
reg  [8:0] _d_uartInBufferNext;
reg  [8:0] _q_uartInBufferNext;
reg  [8:0] _d_uartInBufferTop;
reg  [8:0] _q_uartInBufferTop;
reg  [0:0] _d_uartOutBuffer_wenable0;
reg  [0:0] _q_uartOutBuffer_wenable0;
reg  [8:0] _d_uartOutBuffer_addr0;
reg  [8:0] _q_uartOutBuffer_addr0;
reg  [0:0] _d_uartOutBuffer_wenable1;
reg  [0:0] _q_uartOutBuffer_wenable1;
reg  [7:0] _d_uartOutBuffer_wdata1;
reg  [7:0] _q_uartOutBuffer_wdata1;
reg  [8:0] _d_uartOutBuffer_addr1;
reg  [8:0] _q_uartOutBuffer_addr1;
reg  [8:0] _d_uartOutBufferNext;
reg  [8:0] _q_uartOutBufferNext;
reg  [8:0] _d_uartOutBufferTop;
reg  [8:0] _q_uartOutBufferTop;
reg  [8:0] _d_newuartOutBufferTop;
reg  [8:0] _q_newuartOutBufferTop;
reg  [7:0] _d_led,_q_led;
reg  [7:0] _d_uart_tx_data,_q_uart_tx_data;
reg  [0:0] _d_uart_tx_valid,_q_uart_tx_valid;
reg  [2:0] _d_index,_q_index;
assign out_led = _q_led;
assign out_uart_tx_data = _q_uart_tx_data;
assign out_uart_tx_valid = _q_uart_tx_valid;
assign out_done = (_q_index == 7);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_pc <= 0;
_q_dstack_wenable <= 0;
_q_dstack_wdata <= 0;
_q_dstack_addr <= 0;
_q_stackTop <= 0;
_q_dsp <= 0;
_q_rstack_wenable <= 0;
_q_rstack_wdata <= 0;
_q_rstack_addr <= 0;
_q_rsp <= 0;
_q_rom_addr <= 0;
_q_ram_wenable0 <= 0;
_q_ram_wdata0 <= 0;
_q_ram_addr0 <= 0;
_q_ram_wenable1 <= 0;
_q_ram_addr1 <= 0;
_q_CYCLE <= 0;
_q_INIT <= 0;
_q_copyaddress <= 0;
_q_bramREAD <= 0;
_q_uartInBuffer_wenable0 <= 0;
_q_uartInBuffer_addr0 <= 0;
_q_uartInBuffer_wenable1 <= 0;
_q_uartInBuffer_wdata1 <= 0;
_q_uartInBuffer_addr1 <= 0;
_q_uartInBufferNext <= 0;
_q_uartInBufferTop <= 0;
_q_uartOutBuffer_wenable0 <= 0;
_q_uartOutBuffer_addr0 <= 0;
_q_uartOutBuffer_wenable1 <= 0;
_q_uartOutBuffer_wdata1 <= 0;
_q_uartOutBuffer_addr1 <= 0;
_q_uartOutBufferNext <= 0;
_q_uartOutBufferTop <= 0;
_q_newuartOutBufferTop <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_instruction <= _d_instruction;
_q_pc <= _d_pc;
_q_newPC <= _d_newPC;
_q_dstack_wenable <= _d_dstack_wenable;
_q_dstack_wdata <= _d_dstack_wdata;
_q_dstack_addr <= _d_dstack_addr;
_q_stackTop <= _d_stackTop;
_q_dsp <= _d_dsp;
_q_newDSP <= _d_newDSP;
_q_newStackTop <= _d_newStackTop;
_q_rstack_wenable <= _d_rstack_wenable;
_q_rstack_wdata <= _d_rstack_wdata;
_q_rstack_addr <= _d_rstack_addr;
_q_rsp <= _d_rsp;
_q_newRSP <= _d_newRSP;
_q_rstackWData <= _d_rstackWData;
_q_stackNext <= _d_stackNext;
_q_rStackTop <= _d_rStackTop;
_q_memoryInput <= _d_memoryInput;
_q_rom_addr <= _d_rom_addr;
_q_ram_wenable0 <= _d_ram_wenable0;
_q_ram_wdata0 <= _d_ram_wdata0;
_q_ram_addr0 <= _d_ram_addr0;
_q_ram_wenable1 <= _d_ram_wenable1;
_q_ram_addr1 <= _d_ram_addr1;
_q_CYCLE <= _d_CYCLE;
_q_INIT <= _d_INIT;
_q_copyaddress <= _d_copyaddress;
_q_bramREAD <= _d_bramREAD;
_q_uartInBuffer_wenable0 <= _d_uartInBuffer_wenable0;
_q_uartInBuffer_addr0 <= _d_uartInBuffer_addr0;
_q_uartInBuffer_wenable1 <= _d_uartInBuffer_wenable1;
_q_uartInBuffer_wdata1 <= _d_uartInBuffer_wdata1;
_q_uartInBuffer_addr1 <= _d_uartInBuffer_addr1;
_q_uartInBufferNext <= _d_uartInBufferNext;
_q_uartInBufferTop <= _d_uartInBufferTop;
_q_uartOutBuffer_wenable0 <= _d_uartOutBuffer_wenable0;
_q_uartOutBuffer_addr0 <= _d_uartOutBuffer_addr0;
_q_uartOutBuffer_wenable1 <= _d_uartOutBuffer_wenable1;
_q_uartOutBuffer_wdata1 <= _d_uartOutBuffer_wdata1;
_q_uartOutBuffer_addr1 <= _d_uartOutBuffer_addr1;
_q_uartOutBufferNext <= _d_uartOutBufferNext;
_q_uartOutBufferTop <= _d_uartOutBufferTop;
_q_newuartOutBufferTop <= _d_newuartOutBufferTop;
_q_index <= _d_index;
  end
_q_led <= _d_led;
_q_uart_tx_data <= _d_uart_tx_data;
_q_uart_tx_valid <= _d_uart_tx_valid;
end


M_main_mem_dstack __mem__dstack(
.clock(clock),
.in_dstack_wenable(_d_dstack_wenable),
.in_dstack_wdata(_d_dstack_wdata),
.in_dstack_addr(_d_dstack_addr),
.out_dstack_rdata(_w_mem_dstack_rdata)
);
M_main_mem_rstack __mem__rstack(
.clock(clock),
.in_rstack_wenable(_d_rstack_wenable),
.in_rstack_wdata(_d_rstack_wdata),
.in_rstack_addr(_d_rstack_addr),
.out_rstack_rdata(_w_mem_rstack_rdata)
);
M_main_mem_rom __mem__rom(
.clock(clock),
.in_rom_addr(_d_rom_addr),
.out_rom_rdata(_w_mem_rom_rdata)
);
M_main_mem_ram __mem__ram(
.clock0(clock),
.clock1(clock),
.in_ram_wenable0(_d_ram_wenable0),
.in_ram_wdata0(_d_ram_wdata0),
.in_ram_addr0(_d_ram_addr0),
.in_ram_wenable1(_d_ram_wenable1),
.in_ram_wdata1(_c_ram_wdata1),
.in_ram_addr1(_d_ram_addr1),
.out_ram_rdata0(_w_mem_ram_rdata0),
.out_ram_rdata1(_w_mem_ram_rdata1)
);
M_main_mem_uartInBuffer __mem__uartInBuffer(
.clock0(clock),
.clock1(clock),
.in_uartInBuffer_wenable0(_d_uartInBuffer_wenable0),
.in_uartInBuffer_wdata0(_c_uartInBuffer_wdata0),
.in_uartInBuffer_addr0(_d_uartInBuffer_addr0),
.in_uartInBuffer_wenable1(_d_uartInBuffer_wenable1),
.in_uartInBuffer_wdata1(_d_uartInBuffer_wdata1),
.in_uartInBuffer_addr1(_d_uartInBuffer_addr1),
.out_uartInBuffer_rdata0(_w_mem_uartInBuffer_rdata0),
.out_uartInBuffer_rdata1(_w_mem_uartInBuffer_rdata1)
);
M_main_mem_uartOutBuffer __mem__uartOutBuffer(
.clock0(clock),
.clock1(clock),
.in_uartOutBuffer_wenable0(_d_uartOutBuffer_wenable0),
.in_uartOutBuffer_wdata0(_c_uartOutBuffer_wdata0),
.in_uartOutBuffer_addr0(_d_uartOutBuffer_addr0),
.in_uartOutBuffer_wenable1(_d_uartOutBuffer_wenable1),
.in_uartOutBuffer_wdata1(_d_uartOutBuffer_wdata1),
.in_uartOutBuffer_addr1(_d_uartOutBuffer_addr1),
.out_uartOutBuffer_rdata0(_w_mem_uartOutBuffer_rdata0),
.out_uartOutBuffer_rdata1(_w_mem_uartOutBuffer_rdata1)
);

assign _w_pcPlusOne = _d_pc+1;
assign _w_rdelta = {{7{_d_instruction[3+:1]}},_d_instruction[2+:1]};
assign _w_rstackWrite = (_w_is_call|(_w_is_alu&_d_instruction[6+:1]));
assign _w_dstackWrite = (_w_is_lit|(_w_is_alu&_d_instruction[7+:1]));
assign _w_ddelta = {{7{_d_instruction[1+:1]}},_d_instruction[0+:1]};
assign _w_is_call = (_d_instruction[13+:3]==3'b010);
assign _w_is_lit = _d_instruction[15+:1];
assign _w_is_alu = (_d_instruction[13+:3]==3'b011);
assign _w_immediate = (_d_instruction[0+:15]);

always @* begin
_d_instruction = _q_instruction;
_d_pc = _q_pc;
_d_newPC = _q_newPC;
_d_dstack_wenable = _q_dstack_wenable;
_d_dstack_wdata = _q_dstack_wdata;
_d_dstack_addr = _q_dstack_addr;
_d_stackTop = _q_stackTop;
_d_dsp = _q_dsp;
_d_newDSP = _q_newDSP;
_d_newStackTop = _q_newStackTop;
_d_rstack_wenable = _q_rstack_wenable;
_d_rstack_wdata = _q_rstack_wdata;
_d_rstack_addr = _q_rstack_addr;
_d_rsp = _q_rsp;
_d_newRSP = _q_newRSP;
_d_rstackWData = _q_rstackWData;
_d_stackNext = _q_stackNext;
_d_rStackTop = _q_rStackTop;
_d_memoryInput = _q_memoryInput;
_d_rom_addr = _q_rom_addr;
_d_ram_wenable0 = _q_ram_wenable0;
_d_ram_wdata0 = _q_ram_wdata0;
_d_ram_addr0 = _q_ram_addr0;
_d_ram_wenable1 = _q_ram_wenable1;
_d_ram_addr1 = _q_ram_addr1;
_d_CYCLE = _q_CYCLE;
_d_INIT = _q_INIT;
_d_copyaddress = _q_copyaddress;
_d_bramREAD = _q_bramREAD;
_d_uartInBuffer_wenable0 = _q_uartInBuffer_wenable0;
_d_uartInBuffer_addr0 = _q_uartInBuffer_addr0;
_d_uartInBuffer_wenable1 = _q_uartInBuffer_wenable1;
_d_uartInBuffer_wdata1 = _q_uartInBuffer_wdata1;
_d_uartInBuffer_addr1 = _q_uartInBuffer_addr1;
_d_uartInBufferNext = _q_uartInBufferNext;
_d_uartInBufferTop = _q_uartInBufferTop;
_d_uartOutBuffer_wenable0 = _q_uartOutBuffer_wenable0;
_d_uartOutBuffer_addr0 = _q_uartOutBuffer_addr0;
_d_uartOutBuffer_wenable1 = _q_uartOutBuffer_wenable1;
_d_uartOutBuffer_wdata1 = _q_uartOutBuffer_wdata1;
_d_uartOutBuffer_addr1 = _q_uartOutBuffer_addr1;
_d_uartOutBufferNext = _q_uartOutBufferNext;
_d_uartOutBufferTop = _q_uartOutBufferTop;
_d_newuartOutBufferTop = _q_newuartOutBufferTop;
_d_led = _q_led;
_d_uart_tx_data = _q_uart_tx_data;
_d_uart_tx_valid = _q_uart_tx_valid;
_d_index = _q_index;
// _always_pre
_d_dstack_wenable = 0;
_d_rstack_wenable = 0;
_d_uartInBuffer_wenable0 = 0;
_d_uartInBuffer_wenable1 = 1;
_d_uartInBuffer_addr0 = _q_uartInBufferNext;
_d_uartInBuffer_addr1 = _q_uartInBufferTop;
_d_uartOutBuffer_wenable0 = 0;
_d_uartOutBuffer_wenable1 = 1;
_d_uartOutBuffer_addr0 = _q_uartOutBufferNext;
_d_uartOutBuffer_addr1 = _q_uartOutBufferTop;
_d_index = 7;
case (_q_index)
0: begin
// _top
// var inits
_d_pc = 0;
_d_dstack_wenable = 0;
_d_dstack_wdata = 0;
_d_dstack_addr = 0;
_d_stackTop = 0;
_d_dsp = 0;
_d_rstack_wenable = 0;
_d_rstack_wdata = 0;
_d_rstack_addr = 0;
_d_rsp = 0;
_d_rom_addr = 0;
_d_ram_wenable0 = 0;
_d_ram_wdata0 = 0;
_d_ram_addr0 = 0;
_d_ram_wenable1 = 0;
_d_ram_addr1 = 0;
_d_CYCLE = 0;
_d_INIT = 0;
_d_copyaddress = 0;
_d_bramREAD = 0;
_d_uartInBuffer_wenable0 = 0;
_d_uartInBuffer_addr0 = 0;
_d_uartInBuffer_wenable1 = 0;
_d_uartInBuffer_wdata1 = 0;
_d_uartInBuffer_addr1 = 0;
_d_uartInBufferNext = 0;
_d_uartInBufferTop = 0;
_d_uartOutBuffer_wenable0 = 0;
_d_uartOutBuffer_addr0 = 0;
_d_uartOutBuffer_wenable1 = 0;
_d_uartOutBuffer_wdata1 = 0;
_d_uartOutBuffer_addr1 = 0;
_d_uartOutBufferNext = 0;
_d_uartOutBufferTop = 0;
_d_newuartOutBufferTop = 0;
// --
_d_index = 1;
end
1: begin
// __while__block_1
if (_q_INIT==0) begin
// __block_2
// __block_4
  case (_q_CYCLE)
  0: begin
// __block_6_case
// __block_7
_d_ram_addr0 = _q_copyaddress;
_d_ram_wdata0 = 0;
_d_ram_wenable0 = 1;
// __block_8
  end
  3: begin
// __block_9_case
// __block_10
_d_copyaddress = _q_copyaddress+1;
_d_ram_wenable0 = 0;
// __block_11
  end
  15: begin
// __block_12_case
// __block_13
if (_q_copyaddress==32768) begin
// __block_14
// __block_16
_d_INIT = 1;
_d_copyaddress = 0;
// __block_17
end else begin
// __block_15
end
// __block_18
// __block_19
  end
  default: begin
// __block_20_case
// __block_21
// __block_22
  end
endcase
// __block_5
_d_CYCLE = (_q_CYCLE==15)?0:_q_CYCLE+1;
// __block_23
_d_index = 1;
end else begin
_d_index = 3;
end
end
3: begin
// __while__block_24
if (_q_INIT==1) begin
// __block_25
// __block_27
  case (_q_CYCLE)
  0: begin
// __block_29_case
// __block_30
_d_rom_addr = _q_copyaddress;
// __block_31
  end
  1: begin
// __block_32_case
// __block_33
_d_bramREAD = _w_mem_rom_rdata;
// __block_34
  end
  2: begin
// __block_35_case
// __block_36
_d_ram_addr0 = _q_copyaddress;
_d_ram_wdata0 = _q_bramREAD;
_d_ram_wenable0 = 1;
// __block_37
  end
  14: begin
// __block_38_case
// __block_39
_d_copyaddress = _q_copyaddress+1;
_d_ram_wenable0 = 0;
// __block_40
  end
  15: begin
// __block_41_case
// __block_42
if (_q_copyaddress==4096) begin
// __block_43
// __block_45
_d_INIT = 3;
_d_copyaddress = 0;
// __block_46
end else begin
// __block_44
end
// __block_47
// __block_48
  end
  default: begin
// __block_49_case
// __block_50
// __block_51
  end
endcase
// __block_28
_d_CYCLE = (_q_CYCLE==15)?0:_q_CYCLE+1;
// __block_52
_d_index = 3;
end else begin
_d_index = 5;
end
end
5: begin
// __while__block_53
if (_q_INIT==3) begin
// __block_54
// __block_56
_d_led = _q_instruction;
if (in_uart_rx_valid) begin
// __block_57
// __block_59
_d_uartInBuffer_wdata1 = in_uart_rx_data;
_d_uartInBufferTop = _q_uartInBufferTop+1;
// __block_60
end else begin
// __block_58
end
// __block_61
if (~(_q_uartOutBufferNext==_q_uartOutBufferTop)&~(in_uart_tx_busy)) begin
// __block_62
// __block_64
_d_uart_tx_data = _w_mem_uartOutBuffer_rdata0;
_d_uart_tx_valid = 1;
_d_uartOutBufferNext = _q_uartOutBufferNext+1;
// __block_65
end else begin
// __block_63
end
// __block_66
_d_uartOutBufferTop = _q_newuartOutBufferTop;
  case (_q_CYCLE)
  0: begin
// __block_68_case
// __block_69
_d_stackNext = _w_mem_dstack_rdata;
_d_rStackTop = _w_mem_rstack_rdata;
_d_ram_addr0 = _q_stackTop>>1;
_d_ram_wenable0 = 0;
_d_ram_addr1 = _q_pc;
_d_ram_wenable1 = 0;
// __block_70
  end
  1: begin
// __block_71_case
// __block_72
_d_memoryInput = _w_mem_ram_rdata0;
_d_instruction = _w_mem_ram_rdata1;
// __block_73
  end
  8: begin
// __block_74_case
// __block_75
if (_w_is_lit) begin
// __block_76
// __block_78
_d_newStackTop = _w_immediate;
_d_newPC = _w_pcPlusOne;
_d_newDSP = _q_dsp+1;
_d_newRSP = _q_rsp;
// __block_79
end else begin
// __block_77
// __block_80
  case (_q_instruction[13+:2])
  2'b00: begin
// __block_82_case
// __block_83
_d_newStackTop = _q_stackTop;
_d_newPC = _q_instruction[0+:13];
_d_newDSP = _q_dsp;
_d_newRSP = _q_rsp;
// __block_84
  end
  2'b01: begin
// __block_85_case
// __block_86
_d_newStackTop = _q_stackNext;
_d_newPC = (_q_stackTop==0)?_q_instruction[0+:13]:_w_pcPlusOne;
_d_newDSP = _q_dsp-1;
_d_newRSP = _q_rsp;
// __block_87
  end
  2'b10: begin
// __block_88_case
// __block_89
_d_newStackTop = _q_stackTop;
_d_newPC = _q_instruction[0+:13];
_d_newDSP = _q_dsp;
_d_newRSP = _q_rsp+1;
_d_rstackWData = _w_pcPlusOne<<1;
// __block_90
  end
  2'b11: begin
// __block_91_case
// __block_92
  case (_q_instruction[4+:1])
  1'b0: begin
// __block_94_case
// __block_95
  case (_q_instruction[8+:4])
  4'b0000: begin
// __block_97_case
// __block_98
_d_newStackTop = _q_stackTop;
// __block_99
  end
  4'b0001: begin
// __block_100_case
// __block_101
_d_newStackTop = _q_stackNext;
// __block_102
  end
  4'b0010: begin
// __block_103_case
// __block_104
_d_newStackTop = _q_stackTop+_q_stackNext;
// __block_105
  end
  4'b0011: begin
// __block_106_case
// __block_107
_d_newStackTop = _q_stackTop&_q_stackNext;
// __block_108
  end
  4'b0100: begin
// __block_109_case
// __block_110
_d_newStackTop = _q_stackTop|_q_stackNext;
// __block_111
  end
  4'b0101: begin
// __block_112_case
// __block_113
_d_newStackTop = _q_stackTop^_q_stackNext;
// __block_114
  end
  4'b0110: begin
// __block_115_case
// __block_116
_d_newStackTop = ~_q_stackTop;
// __block_117
  end
  4'b0111: begin
// __block_118_case
// __block_119
_d_newStackTop = {16{(_q_stackNext==_q_stackTop)}};
// __block_120
  end
  4'b1000: begin
// __block_121_case
// __block_122
_d_newStackTop = {16{($signed(_q_stackNext)<$signed(_q_stackTop))}};
// __block_123
  end
  4'b1001: begin
// __block_124_case
// __block_125
_d_newStackTop = _q_stackNext>>_q_stackTop[0+:4];
// __block_126
  end
  4'b1010: begin
// __block_127_case
// __block_128
_d_newStackTop = _q_stackTop-1;
// __block_129
  end
  4'b1011: begin
// __block_130_case
// __block_131
_d_newStackTop = _q_rStackTop;
// __block_132
  end
  4'b1100: begin
// __block_133_case
// __block_134
  case (_q_stackTop)
  16'hf000: begin
// __block_136_case
// __block_137
_d_newStackTop = {8'b0,_w_mem_uartInBuffer_rdata0};
_d_uartInBufferNext = _q_uartInBufferNext+1;
// __block_138
  end
  16'hf001: begin
// __block_139_case
// __block_140
_d_newStackTop = {14'b0,_d_uart_tx_valid,~(_q_uartInBufferNext==_d_uartInBufferTop)};
// __block_141
  end
  16'hf002: begin
// __block_142_case
// __block_143
_d_newStackTop = _d_led;
// __block_144
  end
  16'hf003: begin
// __block_145_case
// __block_146
_d_newStackTop = {12'b0,in_buttons};
// __block_147
  end
  16'hf004: begin
// __block_148_case
// __block_149
_d_newStackTop = in_timer1hz;
// __block_150
  end
  default: begin
// __block_151_case
// __block_152
_d_newStackTop = _q_memoryInput;
// __block_153
  end
endcase
// __block_135
// __block_154
  end
  4'b1101: begin
// __block_155_case
// __block_156
_d_newStackTop = _q_stackNext<<_q_stackTop[0+:4];
// __block_157
  end
  4'b1110: begin
// __block_158_case
// __block_159
_d_newStackTop = {_q_rsp,_q_dsp};
// __block_160
  end
  4'b1111: begin
// __block_161_case
// __block_162
_d_newStackTop = {16{($unsigned(_q_stackNext)<$unsigned(_q_stackTop))}};
// __block_163
  end
endcase
// __block_96
// __block_164
  end
  1'b1: begin
// __block_165_case
// __block_166
  case (_q_instruction[8+:4])
  4'b0000: begin
// __block_168_case
// __block_169
_d_newStackTop = {16{(_q_stackTop==0)}};
// __block_170
  end
  4'b0001: begin
// __block_171_case
// __block_172
_d_newStackTop = ~{16{(_q_stackTop==0)}};
// __block_173
  end
  4'b0010: begin
// __block_174_case
// __block_175
_d_newStackTop = ~{16{(_q_stackNext==_q_stackTop)}};
// __block_176
  end
  4'b0011: begin
// __block_177_case
// __block_178
_d_newStackTop = _q_stackTop+1;
// __block_179
  end
  4'b0100: begin
// __block_180_case
// __block_181
_d_newStackTop = _q_stackTop<<1;
// __block_182
  end
  4'b0101: begin
// __block_183_case
// __block_184
_d_newStackTop = _q_stackTop>>1;
// __block_185
  end
  4'b0110: begin
// __block_186_case
// __block_187
_d_newStackTop = {16{($signed(_q_stackNext)>$signed(_q_stackTop))}};
// __block_188
  end
  4'b0111: begin
// __block_189_case
// __block_190
_d_newStackTop = {16{($unsigned(_q_stackNext)>$unsigned(_q_stackTop))}};
// __block_191
  end
  4'b1000: begin
// __block_192_case
// __block_193
_d_newStackTop = {16{($signed(_q_stackTop)<$signed(0))}};
// __block_194
  end
  4'b1001: begin
// __block_195_case
// __block_196
_d_newStackTop = {16{($signed(_q_stackTop)>$signed(0))}};
// __block_197
  end
  4'b1010: begin
// __block_198_case
// __block_199
_d_newStackTop = ($signed(_q_stackTop)<$signed(0))?-_q_stackTop:_q_stackTop;
// __block_200
  end
  4'b1011: begin
// __block_201_case
// __block_202
_d_newStackTop = ($signed(_q_stackNext)>$signed(_q_stackTop))?_q_stackNext:_q_stackTop;
// __block_203
  end
  4'b1100: begin
// __block_204_case
// __block_205
_d_newStackTop = ($signed(_q_stackNext)<$signed(_q_stackTop))?_q_stackNext:_q_stackTop;
// __block_206
  end
  4'b1101: begin
// __block_207_case
// __block_208
_d_newStackTop = -_q_stackTop;
// __block_209
  end
  4'b1110: begin
// __block_210_case
// __block_211
_d_newStackTop = _q_stackNext-_q_stackTop;
// __block_212
  end
  4'b1111: begin
// __block_213_case
// __block_214
_d_newStackTop = {16{($signed(_q_stackNext)>=$signed(_q_stackTop))}};
// __block_215
  end
endcase
// __block_167
// __block_216
  end
endcase
// __block_93
_d_newDSP = _q_dsp+_w_ddelta;
_d_newRSP = _q_rsp+_w_rdelta;
_d_rstackWData = _q_stackTop;
_d_newPC = (_q_instruction[12+:1])?_q_rStackTop>>1:_w_pcPlusOne;
if (_q_instruction[5+:1]) begin
// __block_217
// __block_219
  case (_q_stackTop)
  default: begin
// __block_221_case
// __block_222
_d_ram_addr0 = _q_stackTop>>1;
_d_ram_wdata0 = _q_stackNext;
_d_ram_wenable0 = 1;
// __block_223
  end
  16'hf000: begin
// __block_224_case
// __block_225
_d_uartOutBuffer_wdata1 = _q_stackNext[0+:8];
_d_newuartOutBufferTop = _d_uartOutBufferTop+1;
// __block_226
  end
  16'hf002: begin
// __block_227_case
// __block_228
_d_led = _q_stackNext;
// __block_229
  end
endcase
// __block_220
// __block_230
end else begin
// __block_218
end
// __block_231
// __block_232
  end
endcase
// __block_81
// __block_233
end
// __block_234
// __block_235
  end
  9: begin
// __block_236_case
// __block_237
if (_w_dstackWrite) begin
// __block_238
// __block_240
_d_dstack_wenable = 1;
_d_dstack_addr = _q_newDSP;
_d_dstack_wdata = _q_stackTop;
// __block_241
end else begin
// __block_239
end
// __block_242
if (_w_rstackWrite) begin
// __block_243
// __block_245
_d_rstack_wenable = 1;
_d_rstack_addr = _q_newRSP;
_d_rstack_wdata = _q_rstackWData;
// __block_246
end else begin
// __block_244
end
// __block_247
// __block_248
  end
  10: begin
// __block_249_case
// __block_250
_d_dsp = _q_newDSP;
_d_pc = _q_newPC;
_d_stackTop = _q_newStackTop;
_d_rsp = _q_newRSP;
_d_dstack_addr = _q_newDSP;
_d_rstack_addr = _q_newRSP;
// __block_251
  end
  12: begin
// __block_252_case
// __block_253
_d_ram_wenable0 = 0;
// __block_254
  end
  default: begin
// __block_255_case
// __block_256
// __block_257
  end
endcase
// __block_67
if (~in_uart_tx_busy&_d_uart_tx_valid) begin
// __block_258
// __block_260
_d_uart_tx_valid = 0;
// __block_261
end else begin
// __block_259
end
// __block_262
_d_CYCLE = _q_CYCLE+1;
// __block_263
_d_index = 5;
end else begin
_d_index = 6;
end
end
6: begin
// __block_55
_d_index = 7;
end
7: begin // end of main
end
default: begin 
_d_index = 7;
 end
endcase
end
endmodule

