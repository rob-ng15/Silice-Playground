`define DE10NANO 1

module SdramVga(
    input clk,
    output reg[7:0] led,

    // SDRAM
    output reg SDRAM_CLK,
    output reg SDRAM_CKE,
    output reg SDRAM_DQML,
    output reg SDRAM_DQMH,
    output reg SDRAM_nCS,
    output reg SDRAM_nWE,
    output reg SDRAM_nCAS,
    output reg SDRAM_nRAS,
    output reg [1:0] SDRAM_BA,
    output reg [12:0] SDRAM_A,
    // inout [15:0] SDRAM_DQ,
    inout [7:0] SDRAM_DQ,

    // VGA
    output reg vga_hs,
    output reg vga_vs,
    output reg [5:0] vga_r,
    output reg [5:0] vga_g,
    output reg [5:0] vga_b,

    // uart via GPIO pins
    output tx,
    input rx,
    
    // user button and switches
    input   BUTTON0,
    input   BUTTON1,
    input   SWITCH0,
    input   SWITCH1,
    input   SWITCH2,
    input   SWITCH3    
);

wire [7:0]  __main_out_led;

wire        __main_out_sdram_clk;
wire        __main_out_sdram_cle;
wire        __main_out_sdram_dqm;
wire        __main_out_sdram_cs;
wire        __main_out_sdram_we;
wire        __main_out_sdram_cas;
wire        __main_out_sdram_ras;
wire [1:0]  __main_out_sdram_ba;
wire [12:0] __main_out_sdram_a;
  
wire        __main_out_vga_hs;
wire        __main_out_vga_vs;
wire [5:0]  __main_out_vga_r;
wire [5:0]  __main_out_vga_g;
wire [5:0]  __main_out_vga_b;

reg [31:0] RST_d;
reg [31:0] RST_q;

reg ready = 0;

always @* begin
  RST_d = RST_q >> 1;
end

always @(posedge clk) begin
  if (ready) begin
    RST_q <= RST_d;
  end else begin
    ready <= 1;
    RST_q <= 32'b111111111111111111111111111111;
  end
end

wire reset_main;
assign reset_main = RST_q[0];
wire run_main;
assign run_main = 1'b1;

// Create 1hz (1 second counter)
reg [31:0] counter50mhz;
reg [15:0] counter1hz;
always @(posedge clk) begin
    if( counter50mhz == 50000000 ) begin
        counter1hz <= counter1hz + 1;
        counter50mhz <= 0;
    end else begin
        counter50mhz <= counter50mhz + 1;
    end
end 

// UART tx and rx
wire [7:0] uart_tx_data;
wire uart_tx_valid;
wire uart_tx_busy;
wire uart_tx_done;
wire [7:0] uart_rx_data;
wire uart_rx_valid;
wire uart_rx_ready;

// UART from https://github.com/jamieiles/uart
uart uart0(
    .din( uart_tx_data ),
    .wr_en( uart_tx_valid ),
    .clk_50m( clk ),
    .tx( tx ),
    .tx_busy( uart_tx_busy ),
    .rx( rx ),
    .rdy( uart_rx_valid ),
    .rdy_clr( uart_rx_ready ),
    .dout( uart_rx_data )
);

// UART from https://github.com/cyrozap/osdvu
//uart uart0(
//    .clk(clk), // The master clock for this module
//    .rst(reset_main), // Synchronous reset
//    .rx(rx), // Incoming serial line
//    .tx(tx), // Outgoing serial line
//    .transmit(uart_tx_valid), // Signal to transmit
//    .tx_byte(uart_tx_data), // Byte to transmit
//    .received(uart_rx_valid), // Indicated that a byte has been received
//    .rx_byte(uart_rx_data), // Byte received
//    .is_receiving(), // Low when receive line is idle
//    .is_transmitting(uart_tx_busy),// Low when transmit line is idle
//    .recv_error() // Indicates error in receiving packet.
//);

M_main __main(
  // CLK and RESET
  .clock(clk),
  .reset(reset_main),
  .in_run(run_main),
  
  // LEDS
  .out_led(__main_out_led),

  // BUTTONS and SWITCHES (combined)
  .in_buttons( {2'b0, SWITCH3, SWITCH2, SWITCH1, SWITCH0, BUTTON1, BUTTON0} ),
  
  .inout_sdram_dq(SDRAM_DQ[7:0]),
  .out_sdram_clk(__main_out_sdram_clk),
  .out_sdram_cle(__main_out_sdram_cle),
  .out_sdram_dqm(__main_out_sdram_dqm),
  .out_sdram_cs(__main_out_sdram_cs),
  .out_sdram_we(__main_out_sdram_we),
  .out_sdram_cas(__main_out_sdram_cas),
  .out_sdram_ras(__main_out_sdram_ras),
  .out_sdram_ba(__main_out_sdram_ba),
  .out_sdram_a(__main_out_sdram_a),
  .out_video_hs(__main_out_vga_hs),
  .out_video_vs(__main_out_vga_vs),
  .out_video_r(__main_out_vga_r),
  .out_video_g(__main_out_vga_g),
  .out_video_b(__main_out_vga_b),

  // UART
  .out_uart_tx_data( uart_tx_data ),
  .out_uart_tx_valid( uart_tx_valid ),
  .in_uart_tx_busy( uart_tx_busy ),
  .in_uart_tx_done( uart_tx_done ),

  .in_uart_rx_data( uart_rx_data ),
  .in_uart_rx_valid( uart_rx_valid ),
  .out_uart_rx_ready( uart_rx_ready ),  
  .in_timer1hz ( counter1hz )
);

always @* begin

  led          = __main_out_led;

  SDRAM_CLK    = __main_out_sdram_clk;
  SDRAM_CKE    = __main_out_sdram_cle;
  SDRAM_DQML   = __main_out_sdram_dqm;
  SDRAM_DQMH   = 0;
  SDRAM_nCS    = __main_out_sdram_cs;
  SDRAM_nWE    = __main_out_sdram_we;
  SDRAM_nCAS   = __main_out_sdram_cas;
  SDRAM_nRAS   = __main_out_sdram_ras;
  SDRAM_BA     = __main_out_sdram_ba;
  SDRAM_A      = __main_out_sdram_a;
  vga_hs       = __main_out_vga_hs;
  vga_vs       = __main_out_vga_vs;
  vga_r        = __main_out_vga_r;
  vga_g        = __main_out_vga_g;
  vga_b        = __main_out_vga_b;

end

endmodule

`timescale 1ns/10ps

module  de10nano_clk_100_25(
	// interface 'refclk'
	input refclk,
	// interface 'reset'
	input rst,
	// interface 'outclk0'
	output outclk_0,
	// interface 'outclk1'
	output outclk_1,
	// interface 'locked'
	output locked
);

	altera_pll #(
		.fractional_vco_multiplier("true"),
		.reference_clock_frequency("50.0 MHz"),
		.operation_mode("direct"),
		.number_of_clocks(2),
		.output_clock_frequency0("100.000000 MHz"),
		.phase_shift0("0 ps"),
		.duty_cycle0(50),
		.output_clock_frequency1("25.000000 MHz"),
		.phase_shift1("0 ps"),
		.duty_cycle1(50),
		.output_clock_frequency2("0 MHz"),
		.phase_shift2("0 ps"),
		.duty_cycle2(50),
		.output_clock_frequency3("0 MHz"),
		.phase_shift3("0 ps"),
		.duty_cycle3(50),
		.output_clock_frequency4("0 MHz"),
		.phase_shift4("0 ps"),
		.duty_cycle4(50),
		.output_clock_frequency5("0 MHz"),
		.phase_shift5("0 ps"),
		.duty_cycle5(50),
		.output_clock_frequency6("0 MHz"),
		.phase_shift6("0 ps"),
		.duty_cycle6(50),
		.output_clock_frequency7("0 MHz"),
		.phase_shift7("0 ps"),
		.duty_cycle7(50),
		.output_clock_frequency8("0 MHz"),
		.phase_shift8("0 ps"),
		.duty_cycle8(50),
		.output_clock_frequency9("0 MHz"),
		.phase_shift9("0 ps"),
		.duty_cycle9(50),
		.output_clock_frequency10("0 MHz"),
		.phase_shift10("0 ps"),
		.duty_cycle10(50),
		.output_clock_frequency11("0 MHz"),
		.phase_shift11("0 ps"),
		.duty_cycle11(50),
		.output_clock_frequency12("0 MHz"),
		.phase_shift12("0 ps"),
		.duty_cycle12(50),
		.output_clock_frequency13("0 MHz"),
		.phase_shift13("0 ps"),
		.duty_cycle13(50),
		.output_clock_frequency14("0 MHz"),
		.phase_shift14("0 ps"),
		.duty_cycle14(50),
		.output_clock_frequency15("0 MHz"),
		.phase_shift15("0 ps"),
		.duty_cycle15(50),
		.output_clock_frequency16("0 MHz"),
		.phase_shift16("0 ps"),
		.duty_cycle16(50),
		.output_clock_frequency17("0 MHz"),
		.phase_shift17("0 ps"),
		.duty_cycle17(50),
		.pll_type("General"),
		.pll_subtype("General")
	) altera_pll_i (
		.rst	(rst),
		.outclk	({outclk_1, outclk_0}),
		.locked	(locked),
		.fboutclk	( ),
		.fbclk	(1'b0),
		.refclk	(refclk)
	);
endmodule



module reset_conditioner (
    input rcclk,
    input in,
    output reg out
  );  
  reg [7:0] counter_d,counter_q;
  always @* begin
    counter_d = counter_q;
    if (counter_q == 0) begin
      out = 0;
    end else begin
      out = 1;
      counter_d = counter_q + 1;
    end
  end  
  always @(posedge rcclk) begin
    if (in == 1'b1) begin
      counter_q <= 1;
    end else begin
      counter_q <= counter_d;
    end
  end 
endmodule


module M_vga (
out_vga_hs,
out_vga_vs,
out_active,
out_vblank,
out_vga_x,
out_vga_y,
in_run,
out_done,
reset,
clock
);
output  [0:0] out_vga_hs;
output  [0:0] out_vga_vs;
output  [0:0] out_active;
output  [0:0] out_vblank;
output  [9:0] out_vga_x;
output  [9:0] out_vga_y;
input in_run;
output out_done;
input reset;
input clock;
wire  [9:0] _c_H_FRT_PORCH;
assign _c_H_FRT_PORCH = 16;
wire  [9:0] _c_H_SYNCH;
assign _c_H_SYNCH = 96;
wire  [9:0] _c_H_BCK_PORCH;
assign _c_H_BCK_PORCH = 48;
wire  [9:0] _c_H_RES;
assign _c_H_RES = 640;
wire  [9:0] _c_V_FRT_PORCH;
assign _c_V_FRT_PORCH = 10;
wire  [9:0] _c_V_SYNCH;
assign _c_V_SYNCH = 2;
wire  [9:0] _c_V_BCK_PORCH;
assign _c_V_BCK_PORCH = 33;
wire  [9:0] _c_V_RES;
assign _c_V_RES = 480;
reg  [9:0] _t_HS_START;
reg  [9:0] _t_HS_END;
reg  [9:0] _t_HA_START;
reg  [9:0] _t_H_END;
reg  [9:0] _t_VS_START;
reg  [9:0] _t_VS_END;
reg  [9:0] _t_VA_START;
reg  [9:0] _t_V_END;

reg  [9:0] _d_xcount;
reg  [9:0] _q_xcount;
reg  [9:0] _d_ycount;
reg  [9:0] _q_ycount;
reg  [0:0] _d_vga_hs,_q_vga_hs;
reg  [0:0] _d_vga_vs,_q_vga_vs;
reg  [0:0] _d_active,_q_active;
reg  [0:0] _d_vblank,_q_vblank;
reg  [9:0] _d_vga_x,_q_vga_x;
reg  [9:0] _d_vga_y,_q_vga_y;
reg  [1:0] _d_index,_q_index;
assign out_vga_hs = _d_vga_hs;
assign out_vga_vs = _d_vga_vs;
assign out_active = _d_active;
assign out_vblank = _d_vblank;
assign out_vga_x = _d_vga_x;
assign out_vga_y = _d_vga_y;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_xcount <= 0;
_q_ycount <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_xcount <= _d_xcount;
_q_ycount <= _d_ycount;
_q_index <= _d_index;
  end
_q_vga_hs <= _d_vga_hs;
_q_vga_vs <= _d_vga_vs;
_q_active <= _d_active;
_q_vblank <= _d_vblank;
_q_vga_x <= _d_vga_x;
_q_vga_y <= _d_vga_y;
end




always @* begin
_d_xcount = _q_xcount;
_d_ycount = _q_ycount;
_d_vga_hs = _q_vga_hs;
_d_vga_vs = _q_vga_vs;
_d_active = _q_active;
_d_vblank = _q_vblank;
_d_vga_x = _q_vga_x;
_d_vga_y = _q_vga_y;
_d_index = _q_index;
_t_HS_START = 0;
_t_HS_END = 0;
_t_HA_START = 0;
_t_H_END = 0;
_t_VS_START = 0;
_t_VS_END = 0;
_t_VA_START = 0;
_t_V_END = 0;
// _always_pre
_t_HS_START = _c_H_FRT_PORCH;
_t_HS_END = _c_H_FRT_PORCH+_c_H_SYNCH;
_t_HA_START = _c_H_FRT_PORCH+_c_H_SYNCH+_c_H_BCK_PORCH;
_t_H_END = _c_H_FRT_PORCH+_c_H_SYNCH+_c_H_BCK_PORCH+_c_H_RES;
_t_VS_START = _c_V_FRT_PORCH;
_t_VS_END = _c_V_FRT_PORCH+_c_V_SYNCH;
_t_VA_START = _c_V_FRT_PORCH+_c_V_SYNCH+_c_V_BCK_PORCH;
_t_V_END = _c_V_FRT_PORCH+_c_V_SYNCH+_c_V_BCK_PORCH+_c_V_RES;
_d_vga_hs = ~((_q_xcount>=_t_HS_START&&_q_xcount<_t_HS_END));
_d_vga_vs = ~((_q_ycount>=_t_VS_START&&_q_ycount<_t_VS_END));
_d_active = (_q_xcount>=_t_HA_START&&_q_xcount<_t_H_END)&&(_q_ycount>=_t_VA_START&&_q_ycount<_t_V_END);
_d_vblank = (_q_ycount<_t_VA_START);
_d_index = 3;
case (_q_index)
0: begin
// _top
// var inits
_t_HS_START = 0;
_t_HS_END = 0;
_t_HA_START = 0;
_t_H_END = 0;
_t_VS_START = 0;
_t_VS_END = 0;
_t_VA_START = 0;
_t_V_END = 0;
_d_xcount = 0;
_d_ycount = 0;
// --
_d_xcount = 0;
_d_ycount = 0;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
if (_d_active) begin
// __block_5
// __block_7
_d_vga_x = _q_xcount-_t_HA_START;
_d_vga_y = _q_ycount-_t_VA_START;
// __block_8
end else begin
// __block_6
end
// __block_9
if (_q_xcount==_t_H_END-1) begin
// __block_10
// __block_12
_d_xcount = 0;
if (_q_ycount==_t_V_END-1) begin
// __block_13
// __block_15
_d_ycount = 0;
// __block_16
end else begin
// __block_14
// __block_17
_d_ycount = _q_ycount+1;
// __block_18
end
// __block_19
// __block_20
end else begin
// __block_11
// __block_21
_d_xcount = _q_xcount+1;
// __block_22
end
// __block_23
// __block_24
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of vga
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_multiplex_display_mem_character(
input      [0:0]             in_character_wenable0,
input       [7:0]     in_character_wdata0,
input      [11:0]                in_character_addr0,
input      [0:0]             in_character_wenable1,
input      [7:0]                 in_character_wdata1,
input      [11:0]                in_character_addr1,
output reg  [7:0]     out_character_rdata0,
output reg  [7:0]     out_character_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2399:0];
always @(posedge clock0) begin
  if (in_character_wenable0) begin
    buffer[in_character_addr0] <= in_character_wdata0;
  end else begin
    out_character_rdata0 <= buffer[in_character_addr0];
  end
end
always @(posedge clock1) begin
  if (in_character_wenable1) begin
    buffer[in_character_addr1] <= in_character_wdata1;
  end else begin
    out_character_rdata1 <= buffer[in_character_addr1];
  end
end

endmodule

module M_multiplex_display_mem_foreground(
input      [0:0]             in_foreground_wenable0,
input       [7:0]     in_foreground_wdata0,
input      [11:0]                in_foreground_addr0,
input      [0:0]             in_foreground_wenable1,
input      [7:0]                 in_foreground_wdata1,
input      [11:0]                in_foreground_addr1,
output reg  [7:0]     out_foreground_rdata0,
output reg  [7:0]     out_foreground_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2399:0];
always @(posedge clock0) begin
  if (in_foreground_wenable0) begin
    buffer[in_foreground_addr0] <= in_foreground_wdata0;
  end else begin
    out_foreground_rdata0 <= buffer[in_foreground_addr0];
  end
end
always @(posedge clock1) begin
  if (in_foreground_wenable1) begin
    buffer[in_foreground_addr1] <= in_foreground_wdata1;
  end else begin
    out_foreground_rdata1 <= buffer[in_foreground_addr1];
  end
end

endmodule

module M_multiplex_display_mem_background(
input      [0:0]             in_background_wenable0,
input       [7:0]     in_background_wdata0,
input      [11:0]                in_background_addr0,
input      [0:0]             in_background_wenable1,
input      [7:0]                 in_background_wdata1,
input      [11:0]                in_background_addr1,
output reg  [7:0]     out_background_rdata0,
output reg  [7:0]     out_background_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[2399:0];
always @(posedge clock0) begin
  if (in_background_wenable0) begin
    buffer[in_background_addr0] <= in_background_wdata0;
  end else begin
    out_background_rdata0 <= buffer[in_background_addr0];
  end
end
always @(posedge clock1) begin
  if (in_background_wenable1) begin
    buffer[in_background_addr1] <= in_background_wdata1;
  end else begin
    out_background_rdata1 <= buffer[in_background_addr1];
  end
end

endmodule

module M_multiplex_display_mem_terminal(
input      [0:0]             in_terminal_wenable0,
input       [7:0]     in_terminal_wdata0,
input      [8:0]                in_terminal_addr0,
input      [0:0]             in_terminal_wenable1,
input      [7:0]                 in_terminal_wdata1,
input      [8:0]                in_terminal_addr1,
output reg  [7:0]     out_terminal_rdata0,
output reg  [7:0]     out_terminal_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[319:0];
always @(posedge clock0) begin
  if (in_terminal_wenable0) begin
    buffer[in_terminal_addr0] <= in_terminal_wdata0;
  end else begin
    out_terminal_rdata0 <= buffer[in_terminal_addr0];
  end
end
always @(posedge clock1) begin
  if (in_terminal_wenable1) begin
    buffer[in_terminal_addr1] <= in_terminal_wdata1;
  end else begin
    out_terminal_rdata1 <= buffer[in_terminal_addr1];
  end
end

endmodule

module M_multiplex_display_mem_bitmap(
input      [0:0]             in_bitmap_wenable0,
input       [7:0]     in_bitmap_wdata0,
input      [18:0]                in_bitmap_addr0,
input      [0:0]             in_bitmap_wenable1,
input      [7:0]                 in_bitmap_wdata1,
input      [18:0]                in_bitmap_addr1,
output reg  [7:0]     out_bitmap_rdata0,
output reg  [7:0]     out_bitmap_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[307199:0];
always @(posedge clock0) begin
  if (in_bitmap_wenable0) begin
    buffer[in_bitmap_addr0] <= in_bitmap_wdata0;
  end else begin
    out_bitmap_rdata0 <= buffer[in_bitmap_addr0];
  end
end
always @(posedge clock1) begin
  if (in_bitmap_wenable1) begin
    buffer[in_bitmap_addr1] <= in_bitmap_wdata1;
  end else begin
    out_bitmap_rdata1 <= buffer[in_bitmap_addr1];
  end
end

endmodule

module M_multiplex_display (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_gpu_x,
in_gpu_y,
in_gpu_param0,
in_gpu_param1,
in_gpu_param2,
in_gpu_param3,
in_gpu_colour,
in_gpu_write,
in_tpu_x,
in_tpu_y,
in_tpu_set,
in_tpu_write,
in_terminal_character,
in_terminal_write,
in_showterminal,
in_showcursor,
in_timer1hz,
out_pix_red,
out_pix_green,
out_pix_blue,
out_gpu_active,
in_run,
out_done,
reset,
clock
);
input  [9:0] in_pix_x;
input  [9:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [9:0] in_gpu_x;
input  [8:0] in_gpu_y;
input  [15:0] in_gpu_param0;
input  [15:0] in_gpu_param1;
input  [15:0] in_gpu_param2;
input  [15:0] in_gpu_param3;
input  [7:0] in_gpu_colour;
input  [1:0] in_gpu_write;
input  [6:0] in_tpu_x;
input  [4:0] in_tpu_y;
input  [7:0] in_tpu_set;
input  [1:0] in_tpu_write;
input  [7:0] in_terminal_character;
input  [0:0] in_terminal_write;
input  [0:0] in_showterminal;
input  [0:0] in_showcursor;
input  [0:0] in_timer1hz;
output  [5:0] out_pix_red;
output  [5:0] out_pix_green;
output  [5:0] out_pix_blue;
output  [7:0] out_gpu_active;
input in_run;
output out_done;
input reset;
input clock;
wire  [7:0] _w_mem_character_rdata0;
wire  [7:0] _w_mem_character_rdata1;
wire  [7:0] _w_mem_foreground_rdata0;
wire  [7:0] _w_mem_foreground_rdata1;
wire  [7:0] _w_mem_background_rdata0;
wire  [7:0] _w_mem_background_rdata1;
wire  [7:0] _w_mem_terminal_rdata0;
wire  [7:0] _w_mem_terminal_rdata1;
wire  [7:0] _w_mem_bitmap_rdata0;
wire  [7:0] _w_mem_bitmap_rdata1;
wire  [7:0] _c_characterGenerator8x16[4095:0];
assign _c_characterGenerator8x16[0] = 8'h00;
assign _c_characterGenerator8x16[1] = 8'h00;
assign _c_characterGenerator8x16[2] = 8'h00;
assign _c_characterGenerator8x16[3] = 8'h00;
assign _c_characterGenerator8x16[4] = 8'h00;
assign _c_characterGenerator8x16[5] = 8'h00;
assign _c_characterGenerator8x16[6] = 8'h00;
assign _c_characterGenerator8x16[7] = 8'h00;
assign _c_characterGenerator8x16[8] = 8'h00;
assign _c_characterGenerator8x16[9] = 8'h00;
assign _c_characterGenerator8x16[10] = 8'h00;
assign _c_characterGenerator8x16[11] = 8'h00;
assign _c_characterGenerator8x16[12] = 8'h00;
assign _c_characterGenerator8x16[13] = 8'h00;
assign _c_characterGenerator8x16[14] = 8'h00;
assign _c_characterGenerator8x16[15] = 8'h00;
assign _c_characterGenerator8x16[16] = 8'h00;
assign _c_characterGenerator8x16[17] = 8'h00;
assign _c_characterGenerator8x16[18] = 8'h7e;
assign _c_characterGenerator8x16[19] = 8'h81;
assign _c_characterGenerator8x16[20] = 8'ha5;
assign _c_characterGenerator8x16[21] = 8'h81;
assign _c_characterGenerator8x16[22] = 8'h81;
assign _c_characterGenerator8x16[23] = 8'hbd;
assign _c_characterGenerator8x16[24] = 8'h99;
assign _c_characterGenerator8x16[25] = 8'h81;
assign _c_characterGenerator8x16[26] = 8'h81;
assign _c_characterGenerator8x16[27] = 8'h7e;
assign _c_characterGenerator8x16[28] = 8'h00;
assign _c_characterGenerator8x16[29] = 8'h00;
assign _c_characterGenerator8x16[30] = 8'h00;
assign _c_characterGenerator8x16[31] = 8'h00;
assign _c_characterGenerator8x16[32] = 8'h00;
assign _c_characterGenerator8x16[33] = 8'h00;
assign _c_characterGenerator8x16[34] = 8'h7e;
assign _c_characterGenerator8x16[35] = 8'hff;
assign _c_characterGenerator8x16[36] = 8'hdb;
assign _c_characterGenerator8x16[37] = 8'hff;
assign _c_characterGenerator8x16[38] = 8'hff;
assign _c_characterGenerator8x16[39] = 8'hc3;
assign _c_characterGenerator8x16[40] = 8'he7;
assign _c_characterGenerator8x16[41] = 8'hff;
assign _c_characterGenerator8x16[42] = 8'hff;
assign _c_characterGenerator8x16[43] = 8'h7e;
assign _c_characterGenerator8x16[44] = 8'h00;
assign _c_characterGenerator8x16[45] = 8'h00;
assign _c_characterGenerator8x16[46] = 8'h00;
assign _c_characterGenerator8x16[47] = 8'h00;
assign _c_characterGenerator8x16[48] = 8'h00;
assign _c_characterGenerator8x16[49] = 8'h00;
assign _c_characterGenerator8x16[50] = 8'h00;
assign _c_characterGenerator8x16[51] = 8'h00;
assign _c_characterGenerator8x16[52] = 8'h6c;
assign _c_characterGenerator8x16[53] = 8'hfe;
assign _c_characterGenerator8x16[54] = 8'hfe;
assign _c_characterGenerator8x16[55] = 8'hfe;
assign _c_characterGenerator8x16[56] = 8'hfe;
assign _c_characterGenerator8x16[57] = 8'h7c;
assign _c_characterGenerator8x16[58] = 8'h38;
assign _c_characterGenerator8x16[59] = 8'h10;
assign _c_characterGenerator8x16[60] = 8'h00;
assign _c_characterGenerator8x16[61] = 8'h00;
assign _c_characterGenerator8x16[62] = 8'h00;
assign _c_characterGenerator8x16[63] = 8'h00;
assign _c_characterGenerator8x16[64] = 8'h00;
assign _c_characterGenerator8x16[65] = 8'h00;
assign _c_characterGenerator8x16[66] = 8'h00;
assign _c_characterGenerator8x16[67] = 8'h00;
assign _c_characterGenerator8x16[68] = 8'h10;
assign _c_characterGenerator8x16[69] = 8'h38;
assign _c_characterGenerator8x16[70] = 8'h7c;
assign _c_characterGenerator8x16[71] = 8'hfe;
assign _c_characterGenerator8x16[72] = 8'h7c;
assign _c_characterGenerator8x16[73] = 8'h38;
assign _c_characterGenerator8x16[74] = 8'h10;
assign _c_characterGenerator8x16[75] = 8'h00;
assign _c_characterGenerator8x16[76] = 8'h00;
assign _c_characterGenerator8x16[77] = 8'h00;
assign _c_characterGenerator8x16[78] = 8'h00;
assign _c_characterGenerator8x16[79] = 8'h00;
assign _c_characterGenerator8x16[80] = 8'h00;
assign _c_characterGenerator8x16[81] = 8'h00;
assign _c_characterGenerator8x16[82] = 8'h00;
assign _c_characterGenerator8x16[83] = 8'h18;
assign _c_characterGenerator8x16[84] = 8'h3c;
assign _c_characterGenerator8x16[85] = 8'h3c;
assign _c_characterGenerator8x16[86] = 8'he7;
assign _c_characterGenerator8x16[87] = 8'he7;
assign _c_characterGenerator8x16[88] = 8'he7;
assign _c_characterGenerator8x16[89] = 8'h18;
assign _c_characterGenerator8x16[90] = 8'h18;
assign _c_characterGenerator8x16[91] = 8'h3c;
assign _c_characterGenerator8x16[92] = 8'h00;
assign _c_characterGenerator8x16[93] = 8'h00;
assign _c_characterGenerator8x16[94] = 8'h00;
assign _c_characterGenerator8x16[95] = 8'h00;
assign _c_characterGenerator8x16[96] = 8'h00;
assign _c_characterGenerator8x16[97] = 8'h00;
assign _c_characterGenerator8x16[98] = 8'h00;
assign _c_characterGenerator8x16[99] = 8'h18;
assign _c_characterGenerator8x16[100] = 8'h3c;
assign _c_characterGenerator8x16[101] = 8'h7e;
assign _c_characterGenerator8x16[102] = 8'hff;
assign _c_characterGenerator8x16[103] = 8'hff;
assign _c_characterGenerator8x16[104] = 8'h7e;
assign _c_characterGenerator8x16[105] = 8'h18;
assign _c_characterGenerator8x16[106] = 8'h18;
assign _c_characterGenerator8x16[107] = 8'h3c;
assign _c_characterGenerator8x16[108] = 8'h00;
assign _c_characterGenerator8x16[109] = 8'h00;
assign _c_characterGenerator8x16[110] = 8'h00;
assign _c_characterGenerator8x16[111] = 8'h00;
assign _c_characterGenerator8x16[112] = 8'h00;
assign _c_characterGenerator8x16[113] = 8'h00;
assign _c_characterGenerator8x16[114] = 8'h00;
assign _c_characterGenerator8x16[115] = 8'h00;
assign _c_characterGenerator8x16[116] = 8'h00;
assign _c_characterGenerator8x16[117] = 8'h00;
assign _c_characterGenerator8x16[118] = 8'h18;
assign _c_characterGenerator8x16[119] = 8'h3c;
assign _c_characterGenerator8x16[120] = 8'h3c;
assign _c_characterGenerator8x16[121] = 8'h18;
assign _c_characterGenerator8x16[122] = 8'h00;
assign _c_characterGenerator8x16[123] = 8'h00;
assign _c_characterGenerator8x16[124] = 8'h00;
assign _c_characterGenerator8x16[125] = 8'h00;
assign _c_characterGenerator8x16[126] = 8'h00;
assign _c_characterGenerator8x16[127] = 8'h00;
assign _c_characterGenerator8x16[128] = 8'hff;
assign _c_characterGenerator8x16[129] = 8'hff;
assign _c_characterGenerator8x16[130] = 8'hff;
assign _c_characterGenerator8x16[131] = 8'hff;
assign _c_characterGenerator8x16[132] = 8'hff;
assign _c_characterGenerator8x16[133] = 8'hff;
assign _c_characterGenerator8x16[134] = 8'he7;
assign _c_characterGenerator8x16[135] = 8'hc3;
assign _c_characterGenerator8x16[136] = 8'hc3;
assign _c_characterGenerator8x16[137] = 8'he7;
assign _c_characterGenerator8x16[138] = 8'hff;
assign _c_characterGenerator8x16[139] = 8'hff;
assign _c_characterGenerator8x16[140] = 8'hff;
assign _c_characterGenerator8x16[141] = 8'hff;
assign _c_characterGenerator8x16[142] = 8'hff;
assign _c_characterGenerator8x16[143] = 8'hff;
assign _c_characterGenerator8x16[144] = 8'h00;
assign _c_characterGenerator8x16[145] = 8'h00;
assign _c_characterGenerator8x16[146] = 8'h00;
assign _c_characterGenerator8x16[147] = 8'h00;
assign _c_characterGenerator8x16[148] = 8'h00;
assign _c_characterGenerator8x16[149] = 8'h3c;
assign _c_characterGenerator8x16[150] = 8'h66;
assign _c_characterGenerator8x16[151] = 8'h42;
assign _c_characterGenerator8x16[152] = 8'h42;
assign _c_characterGenerator8x16[153] = 8'h66;
assign _c_characterGenerator8x16[154] = 8'h3c;
assign _c_characterGenerator8x16[155] = 8'h00;
assign _c_characterGenerator8x16[156] = 8'h00;
assign _c_characterGenerator8x16[157] = 8'h00;
assign _c_characterGenerator8x16[158] = 8'h00;
assign _c_characterGenerator8x16[159] = 8'h00;
assign _c_characterGenerator8x16[160] = 8'hff;
assign _c_characterGenerator8x16[161] = 8'hff;
assign _c_characterGenerator8x16[162] = 8'hff;
assign _c_characterGenerator8x16[163] = 8'hff;
assign _c_characterGenerator8x16[164] = 8'hff;
assign _c_characterGenerator8x16[165] = 8'hc3;
assign _c_characterGenerator8x16[166] = 8'h99;
assign _c_characterGenerator8x16[167] = 8'hbd;
assign _c_characterGenerator8x16[168] = 8'hbd;
assign _c_characterGenerator8x16[169] = 8'h99;
assign _c_characterGenerator8x16[170] = 8'hc3;
assign _c_characterGenerator8x16[171] = 8'hff;
assign _c_characterGenerator8x16[172] = 8'hff;
assign _c_characterGenerator8x16[173] = 8'hff;
assign _c_characterGenerator8x16[174] = 8'hff;
assign _c_characterGenerator8x16[175] = 8'hff;
assign _c_characterGenerator8x16[176] = 8'h00;
assign _c_characterGenerator8x16[177] = 8'h00;
assign _c_characterGenerator8x16[178] = 8'h1e;
assign _c_characterGenerator8x16[179] = 8'h0e;
assign _c_characterGenerator8x16[180] = 8'h1a;
assign _c_characterGenerator8x16[181] = 8'h32;
assign _c_characterGenerator8x16[182] = 8'h78;
assign _c_characterGenerator8x16[183] = 8'hcc;
assign _c_characterGenerator8x16[184] = 8'hcc;
assign _c_characterGenerator8x16[185] = 8'hcc;
assign _c_characterGenerator8x16[186] = 8'hcc;
assign _c_characterGenerator8x16[187] = 8'h78;
assign _c_characterGenerator8x16[188] = 8'h00;
assign _c_characterGenerator8x16[189] = 8'h00;
assign _c_characterGenerator8x16[190] = 8'h00;
assign _c_characterGenerator8x16[191] = 8'h00;
assign _c_characterGenerator8x16[192] = 8'h00;
assign _c_characterGenerator8x16[193] = 8'h00;
assign _c_characterGenerator8x16[194] = 8'h3c;
assign _c_characterGenerator8x16[195] = 8'h66;
assign _c_characterGenerator8x16[196] = 8'h66;
assign _c_characterGenerator8x16[197] = 8'h66;
assign _c_characterGenerator8x16[198] = 8'h66;
assign _c_characterGenerator8x16[199] = 8'h3c;
assign _c_characterGenerator8x16[200] = 8'h18;
assign _c_characterGenerator8x16[201] = 8'h7e;
assign _c_characterGenerator8x16[202] = 8'h18;
assign _c_characterGenerator8x16[203] = 8'h18;
assign _c_characterGenerator8x16[204] = 8'h00;
assign _c_characterGenerator8x16[205] = 8'h00;
assign _c_characterGenerator8x16[206] = 8'h00;
assign _c_characterGenerator8x16[207] = 8'h00;
assign _c_characterGenerator8x16[208] = 8'h00;
assign _c_characterGenerator8x16[209] = 8'h00;
assign _c_characterGenerator8x16[210] = 8'h3f;
assign _c_characterGenerator8x16[211] = 8'h33;
assign _c_characterGenerator8x16[212] = 8'h3f;
assign _c_characterGenerator8x16[213] = 8'h30;
assign _c_characterGenerator8x16[214] = 8'h30;
assign _c_characterGenerator8x16[215] = 8'h30;
assign _c_characterGenerator8x16[216] = 8'h30;
assign _c_characterGenerator8x16[217] = 8'h70;
assign _c_characterGenerator8x16[218] = 8'hf0;
assign _c_characterGenerator8x16[219] = 8'he0;
assign _c_characterGenerator8x16[220] = 8'h00;
assign _c_characterGenerator8x16[221] = 8'h00;
assign _c_characterGenerator8x16[222] = 8'h00;
assign _c_characterGenerator8x16[223] = 8'h00;
assign _c_characterGenerator8x16[224] = 8'h00;
assign _c_characterGenerator8x16[225] = 8'h00;
assign _c_characterGenerator8x16[226] = 8'h7f;
assign _c_characterGenerator8x16[227] = 8'h63;
assign _c_characterGenerator8x16[228] = 8'h7f;
assign _c_characterGenerator8x16[229] = 8'h63;
assign _c_characterGenerator8x16[230] = 8'h63;
assign _c_characterGenerator8x16[231] = 8'h63;
assign _c_characterGenerator8x16[232] = 8'h63;
assign _c_characterGenerator8x16[233] = 8'h67;
assign _c_characterGenerator8x16[234] = 8'he7;
assign _c_characterGenerator8x16[235] = 8'he6;
assign _c_characterGenerator8x16[236] = 8'hc0;
assign _c_characterGenerator8x16[237] = 8'h00;
assign _c_characterGenerator8x16[238] = 8'h00;
assign _c_characterGenerator8x16[239] = 8'h00;
assign _c_characterGenerator8x16[240] = 8'h00;
assign _c_characterGenerator8x16[241] = 8'h00;
assign _c_characterGenerator8x16[242] = 8'h00;
assign _c_characterGenerator8x16[243] = 8'h18;
assign _c_characterGenerator8x16[244] = 8'h18;
assign _c_characterGenerator8x16[245] = 8'hdb;
assign _c_characterGenerator8x16[246] = 8'h3c;
assign _c_characterGenerator8x16[247] = 8'he7;
assign _c_characterGenerator8x16[248] = 8'h3c;
assign _c_characterGenerator8x16[249] = 8'hdb;
assign _c_characterGenerator8x16[250] = 8'h18;
assign _c_characterGenerator8x16[251] = 8'h18;
assign _c_characterGenerator8x16[252] = 8'h00;
assign _c_characterGenerator8x16[253] = 8'h00;
assign _c_characterGenerator8x16[254] = 8'h00;
assign _c_characterGenerator8x16[255] = 8'h00;
assign _c_characterGenerator8x16[256] = 8'h00;
assign _c_characterGenerator8x16[257] = 8'h80;
assign _c_characterGenerator8x16[258] = 8'hc0;
assign _c_characterGenerator8x16[259] = 8'he0;
assign _c_characterGenerator8x16[260] = 8'hf0;
assign _c_characterGenerator8x16[261] = 8'hf8;
assign _c_characterGenerator8x16[262] = 8'hfe;
assign _c_characterGenerator8x16[263] = 8'hf8;
assign _c_characterGenerator8x16[264] = 8'hf0;
assign _c_characterGenerator8x16[265] = 8'he0;
assign _c_characterGenerator8x16[266] = 8'hc0;
assign _c_characterGenerator8x16[267] = 8'h80;
assign _c_characterGenerator8x16[268] = 8'h00;
assign _c_characterGenerator8x16[269] = 8'h00;
assign _c_characterGenerator8x16[270] = 8'h00;
assign _c_characterGenerator8x16[271] = 8'h00;
assign _c_characterGenerator8x16[272] = 8'h00;
assign _c_characterGenerator8x16[273] = 8'h02;
assign _c_characterGenerator8x16[274] = 8'h06;
assign _c_characterGenerator8x16[275] = 8'h0e;
assign _c_characterGenerator8x16[276] = 8'h1e;
assign _c_characterGenerator8x16[277] = 8'h3e;
assign _c_characterGenerator8x16[278] = 8'hfe;
assign _c_characterGenerator8x16[279] = 8'h3e;
assign _c_characterGenerator8x16[280] = 8'h1e;
assign _c_characterGenerator8x16[281] = 8'h0e;
assign _c_characterGenerator8x16[282] = 8'h06;
assign _c_characterGenerator8x16[283] = 8'h02;
assign _c_characterGenerator8x16[284] = 8'h00;
assign _c_characterGenerator8x16[285] = 8'h00;
assign _c_characterGenerator8x16[286] = 8'h00;
assign _c_characterGenerator8x16[287] = 8'h00;
assign _c_characterGenerator8x16[288] = 8'h00;
assign _c_characterGenerator8x16[289] = 8'h00;
assign _c_characterGenerator8x16[290] = 8'h18;
assign _c_characterGenerator8x16[291] = 8'h3c;
assign _c_characterGenerator8x16[292] = 8'h7e;
assign _c_characterGenerator8x16[293] = 8'h18;
assign _c_characterGenerator8x16[294] = 8'h18;
assign _c_characterGenerator8x16[295] = 8'h18;
assign _c_characterGenerator8x16[296] = 8'h7e;
assign _c_characterGenerator8x16[297] = 8'h3c;
assign _c_characterGenerator8x16[298] = 8'h18;
assign _c_characterGenerator8x16[299] = 8'h00;
assign _c_characterGenerator8x16[300] = 8'h00;
assign _c_characterGenerator8x16[301] = 8'h00;
assign _c_characterGenerator8x16[302] = 8'h00;
assign _c_characterGenerator8x16[303] = 8'h00;
assign _c_characterGenerator8x16[304] = 8'h00;
assign _c_characterGenerator8x16[305] = 8'h00;
assign _c_characterGenerator8x16[306] = 8'h66;
assign _c_characterGenerator8x16[307] = 8'h66;
assign _c_characterGenerator8x16[308] = 8'h66;
assign _c_characterGenerator8x16[309] = 8'h66;
assign _c_characterGenerator8x16[310] = 8'h66;
assign _c_characterGenerator8x16[311] = 8'h66;
assign _c_characterGenerator8x16[312] = 8'h66;
assign _c_characterGenerator8x16[313] = 8'h00;
assign _c_characterGenerator8x16[314] = 8'h66;
assign _c_characterGenerator8x16[315] = 8'h66;
assign _c_characterGenerator8x16[316] = 8'h00;
assign _c_characterGenerator8x16[317] = 8'h00;
assign _c_characterGenerator8x16[318] = 8'h00;
assign _c_characterGenerator8x16[319] = 8'h00;
assign _c_characterGenerator8x16[320] = 8'h00;
assign _c_characterGenerator8x16[321] = 8'h00;
assign _c_characterGenerator8x16[322] = 8'h7f;
assign _c_characterGenerator8x16[323] = 8'hdb;
assign _c_characterGenerator8x16[324] = 8'hdb;
assign _c_characterGenerator8x16[325] = 8'hdb;
assign _c_characterGenerator8x16[326] = 8'h7b;
assign _c_characterGenerator8x16[327] = 8'h1b;
assign _c_characterGenerator8x16[328] = 8'h1b;
assign _c_characterGenerator8x16[329] = 8'h1b;
assign _c_characterGenerator8x16[330] = 8'h1b;
assign _c_characterGenerator8x16[331] = 8'h1b;
assign _c_characterGenerator8x16[332] = 8'h00;
assign _c_characterGenerator8x16[333] = 8'h00;
assign _c_characterGenerator8x16[334] = 8'h00;
assign _c_characterGenerator8x16[335] = 8'h00;
assign _c_characterGenerator8x16[336] = 8'h00;
assign _c_characterGenerator8x16[337] = 8'h7c;
assign _c_characterGenerator8x16[338] = 8'hc6;
assign _c_characterGenerator8x16[339] = 8'h60;
assign _c_characterGenerator8x16[340] = 8'h38;
assign _c_characterGenerator8x16[341] = 8'h6c;
assign _c_characterGenerator8x16[342] = 8'hc6;
assign _c_characterGenerator8x16[343] = 8'hc6;
assign _c_characterGenerator8x16[344] = 8'h6c;
assign _c_characterGenerator8x16[345] = 8'h38;
assign _c_characterGenerator8x16[346] = 8'h0c;
assign _c_characterGenerator8x16[347] = 8'hc6;
assign _c_characterGenerator8x16[348] = 8'h7c;
assign _c_characterGenerator8x16[349] = 8'h00;
assign _c_characterGenerator8x16[350] = 8'h00;
assign _c_characterGenerator8x16[351] = 8'h00;
assign _c_characterGenerator8x16[352] = 8'h00;
assign _c_characterGenerator8x16[353] = 8'h00;
assign _c_characterGenerator8x16[354] = 8'h00;
assign _c_characterGenerator8x16[355] = 8'h00;
assign _c_characterGenerator8x16[356] = 8'h00;
assign _c_characterGenerator8x16[357] = 8'h00;
assign _c_characterGenerator8x16[358] = 8'h00;
assign _c_characterGenerator8x16[359] = 8'h00;
assign _c_characterGenerator8x16[360] = 8'hfe;
assign _c_characterGenerator8x16[361] = 8'hfe;
assign _c_characterGenerator8x16[362] = 8'hfe;
assign _c_characterGenerator8x16[363] = 8'hfe;
assign _c_characterGenerator8x16[364] = 8'h00;
assign _c_characterGenerator8x16[365] = 8'h00;
assign _c_characterGenerator8x16[366] = 8'h00;
assign _c_characterGenerator8x16[367] = 8'h00;
assign _c_characterGenerator8x16[368] = 8'h00;
assign _c_characterGenerator8x16[369] = 8'h00;
assign _c_characterGenerator8x16[370] = 8'h18;
assign _c_characterGenerator8x16[371] = 8'h3c;
assign _c_characterGenerator8x16[372] = 8'h7e;
assign _c_characterGenerator8x16[373] = 8'h18;
assign _c_characterGenerator8x16[374] = 8'h18;
assign _c_characterGenerator8x16[375] = 8'h18;
assign _c_characterGenerator8x16[376] = 8'h7e;
assign _c_characterGenerator8x16[377] = 8'h3c;
assign _c_characterGenerator8x16[378] = 8'h18;
assign _c_characterGenerator8x16[379] = 8'h7e;
assign _c_characterGenerator8x16[380] = 8'h00;
assign _c_characterGenerator8x16[381] = 8'h00;
assign _c_characterGenerator8x16[382] = 8'h00;
assign _c_characterGenerator8x16[383] = 8'h00;
assign _c_characterGenerator8x16[384] = 8'h00;
assign _c_characterGenerator8x16[385] = 8'h00;
assign _c_characterGenerator8x16[386] = 8'h18;
assign _c_characterGenerator8x16[387] = 8'h3c;
assign _c_characterGenerator8x16[388] = 8'h7e;
assign _c_characterGenerator8x16[389] = 8'h18;
assign _c_characterGenerator8x16[390] = 8'h18;
assign _c_characterGenerator8x16[391] = 8'h18;
assign _c_characterGenerator8x16[392] = 8'h18;
assign _c_characterGenerator8x16[393] = 8'h18;
assign _c_characterGenerator8x16[394] = 8'h18;
assign _c_characterGenerator8x16[395] = 8'h18;
assign _c_characterGenerator8x16[396] = 8'h00;
assign _c_characterGenerator8x16[397] = 8'h00;
assign _c_characterGenerator8x16[398] = 8'h00;
assign _c_characterGenerator8x16[399] = 8'h00;
assign _c_characterGenerator8x16[400] = 8'h00;
assign _c_characterGenerator8x16[401] = 8'h00;
assign _c_characterGenerator8x16[402] = 8'h18;
assign _c_characterGenerator8x16[403] = 8'h18;
assign _c_characterGenerator8x16[404] = 8'h18;
assign _c_characterGenerator8x16[405] = 8'h18;
assign _c_characterGenerator8x16[406] = 8'h18;
assign _c_characterGenerator8x16[407] = 8'h18;
assign _c_characterGenerator8x16[408] = 8'h18;
assign _c_characterGenerator8x16[409] = 8'h7e;
assign _c_characterGenerator8x16[410] = 8'h3c;
assign _c_characterGenerator8x16[411] = 8'h18;
assign _c_characterGenerator8x16[412] = 8'h00;
assign _c_characterGenerator8x16[413] = 8'h00;
assign _c_characterGenerator8x16[414] = 8'h00;
assign _c_characterGenerator8x16[415] = 8'h00;
assign _c_characterGenerator8x16[416] = 8'h00;
assign _c_characterGenerator8x16[417] = 8'h00;
assign _c_characterGenerator8x16[418] = 8'h00;
assign _c_characterGenerator8x16[419] = 8'h00;
assign _c_characterGenerator8x16[420] = 8'h00;
assign _c_characterGenerator8x16[421] = 8'h18;
assign _c_characterGenerator8x16[422] = 8'h0c;
assign _c_characterGenerator8x16[423] = 8'hfe;
assign _c_characterGenerator8x16[424] = 8'h0c;
assign _c_characterGenerator8x16[425] = 8'h18;
assign _c_characterGenerator8x16[426] = 8'h00;
assign _c_characterGenerator8x16[427] = 8'h00;
assign _c_characterGenerator8x16[428] = 8'h00;
assign _c_characterGenerator8x16[429] = 8'h00;
assign _c_characterGenerator8x16[430] = 8'h00;
assign _c_characterGenerator8x16[431] = 8'h00;
assign _c_characterGenerator8x16[432] = 8'h00;
assign _c_characterGenerator8x16[433] = 8'h00;
assign _c_characterGenerator8x16[434] = 8'h00;
assign _c_characterGenerator8x16[435] = 8'h00;
assign _c_characterGenerator8x16[436] = 8'h00;
assign _c_characterGenerator8x16[437] = 8'h30;
assign _c_characterGenerator8x16[438] = 8'h60;
assign _c_characterGenerator8x16[439] = 8'hfe;
assign _c_characterGenerator8x16[440] = 8'h60;
assign _c_characterGenerator8x16[441] = 8'h30;
assign _c_characterGenerator8x16[442] = 8'h00;
assign _c_characterGenerator8x16[443] = 8'h00;
assign _c_characterGenerator8x16[444] = 8'h00;
assign _c_characterGenerator8x16[445] = 8'h00;
assign _c_characterGenerator8x16[446] = 8'h00;
assign _c_characterGenerator8x16[447] = 8'h00;
assign _c_characterGenerator8x16[448] = 8'h00;
assign _c_characterGenerator8x16[449] = 8'h00;
assign _c_characterGenerator8x16[450] = 8'h00;
assign _c_characterGenerator8x16[451] = 8'h00;
assign _c_characterGenerator8x16[452] = 8'h00;
assign _c_characterGenerator8x16[453] = 8'h00;
assign _c_characterGenerator8x16[454] = 8'hc0;
assign _c_characterGenerator8x16[455] = 8'hc0;
assign _c_characterGenerator8x16[456] = 8'hc0;
assign _c_characterGenerator8x16[457] = 8'hfe;
assign _c_characterGenerator8x16[458] = 8'h00;
assign _c_characterGenerator8x16[459] = 8'h00;
assign _c_characterGenerator8x16[460] = 8'h00;
assign _c_characterGenerator8x16[461] = 8'h00;
assign _c_characterGenerator8x16[462] = 8'h00;
assign _c_characterGenerator8x16[463] = 8'h00;
assign _c_characterGenerator8x16[464] = 8'h00;
assign _c_characterGenerator8x16[465] = 8'h00;
assign _c_characterGenerator8x16[466] = 8'h00;
assign _c_characterGenerator8x16[467] = 8'h00;
assign _c_characterGenerator8x16[468] = 8'h00;
assign _c_characterGenerator8x16[469] = 8'h28;
assign _c_characterGenerator8x16[470] = 8'h6c;
assign _c_characterGenerator8x16[471] = 8'hfe;
assign _c_characterGenerator8x16[472] = 8'h6c;
assign _c_characterGenerator8x16[473] = 8'h28;
assign _c_characterGenerator8x16[474] = 8'h00;
assign _c_characterGenerator8x16[475] = 8'h00;
assign _c_characterGenerator8x16[476] = 8'h00;
assign _c_characterGenerator8x16[477] = 8'h00;
assign _c_characterGenerator8x16[478] = 8'h00;
assign _c_characterGenerator8x16[479] = 8'h00;
assign _c_characterGenerator8x16[480] = 8'h00;
assign _c_characterGenerator8x16[481] = 8'h00;
assign _c_characterGenerator8x16[482] = 8'h00;
assign _c_characterGenerator8x16[483] = 8'h00;
assign _c_characterGenerator8x16[484] = 8'h10;
assign _c_characterGenerator8x16[485] = 8'h38;
assign _c_characterGenerator8x16[486] = 8'h38;
assign _c_characterGenerator8x16[487] = 8'h7c;
assign _c_characterGenerator8x16[488] = 8'h7c;
assign _c_characterGenerator8x16[489] = 8'hfe;
assign _c_characterGenerator8x16[490] = 8'hfe;
assign _c_characterGenerator8x16[491] = 8'h00;
assign _c_characterGenerator8x16[492] = 8'h00;
assign _c_characterGenerator8x16[493] = 8'h00;
assign _c_characterGenerator8x16[494] = 8'h00;
assign _c_characterGenerator8x16[495] = 8'h00;
assign _c_characterGenerator8x16[496] = 8'h00;
assign _c_characterGenerator8x16[497] = 8'h00;
assign _c_characterGenerator8x16[498] = 8'h00;
assign _c_characterGenerator8x16[499] = 8'h00;
assign _c_characterGenerator8x16[500] = 8'hfe;
assign _c_characterGenerator8x16[501] = 8'hfe;
assign _c_characterGenerator8x16[502] = 8'h7c;
assign _c_characterGenerator8x16[503] = 8'h7c;
assign _c_characterGenerator8x16[504] = 8'h38;
assign _c_characterGenerator8x16[505] = 8'h38;
assign _c_characterGenerator8x16[506] = 8'h10;
assign _c_characterGenerator8x16[507] = 8'h00;
assign _c_characterGenerator8x16[508] = 8'h00;
assign _c_characterGenerator8x16[509] = 8'h00;
assign _c_characterGenerator8x16[510] = 8'h00;
assign _c_characterGenerator8x16[511] = 8'h00;
assign _c_characterGenerator8x16[512] = 8'h00;
assign _c_characterGenerator8x16[513] = 8'h00;
assign _c_characterGenerator8x16[514] = 8'h00;
assign _c_characterGenerator8x16[515] = 8'h00;
assign _c_characterGenerator8x16[516] = 8'h00;
assign _c_characterGenerator8x16[517] = 8'h00;
assign _c_characterGenerator8x16[518] = 8'h00;
assign _c_characterGenerator8x16[519] = 8'h00;
assign _c_characterGenerator8x16[520] = 8'h00;
assign _c_characterGenerator8x16[521] = 8'h00;
assign _c_characterGenerator8x16[522] = 8'h00;
assign _c_characterGenerator8x16[523] = 8'h00;
assign _c_characterGenerator8x16[524] = 8'h00;
assign _c_characterGenerator8x16[525] = 8'h00;
assign _c_characterGenerator8x16[526] = 8'h00;
assign _c_characterGenerator8x16[527] = 8'h00;
assign _c_characterGenerator8x16[528] = 8'h00;
assign _c_characterGenerator8x16[529] = 8'h00;
assign _c_characterGenerator8x16[530] = 8'h18;
assign _c_characterGenerator8x16[531] = 8'h3c;
assign _c_characterGenerator8x16[532] = 8'h3c;
assign _c_characterGenerator8x16[533] = 8'h3c;
assign _c_characterGenerator8x16[534] = 8'h18;
assign _c_characterGenerator8x16[535] = 8'h18;
assign _c_characterGenerator8x16[536] = 8'h18;
assign _c_characterGenerator8x16[537] = 8'h00;
assign _c_characterGenerator8x16[538] = 8'h18;
assign _c_characterGenerator8x16[539] = 8'h18;
assign _c_characterGenerator8x16[540] = 8'h00;
assign _c_characterGenerator8x16[541] = 8'h00;
assign _c_characterGenerator8x16[542] = 8'h00;
assign _c_characterGenerator8x16[543] = 8'h00;
assign _c_characterGenerator8x16[544] = 8'h00;
assign _c_characterGenerator8x16[545] = 8'h66;
assign _c_characterGenerator8x16[546] = 8'h66;
assign _c_characterGenerator8x16[547] = 8'h66;
assign _c_characterGenerator8x16[548] = 8'h24;
assign _c_characterGenerator8x16[549] = 8'h00;
assign _c_characterGenerator8x16[550] = 8'h00;
assign _c_characterGenerator8x16[551] = 8'h00;
assign _c_characterGenerator8x16[552] = 8'h00;
assign _c_characterGenerator8x16[553] = 8'h00;
assign _c_characterGenerator8x16[554] = 8'h00;
assign _c_characterGenerator8x16[555] = 8'h00;
assign _c_characterGenerator8x16[556] = 8'h00;
assign _c_characterGenerator8x16[557] = 8'h00;
assign _c_characterGenerator8x16[558] = 8'h00;
assign _c_characterGenerator8x16[559] = 8'h00;
assign _c_characterGenerator8x16[560] = 8'h00;
assign _c_characterGenerator8x16[561] = 8'h00;
assign _c_characterGenerator8x16[562] = 8'h00;
assign _c_characterGenerator8x16[563] = 8'h6c;
assign _c_characterGenerator8x16[564] = 8'h6c;
assign _c_characterGenerator8x16[565] = 8'hfe;
assign _c_characterGenerator8x16[566] = 8'h6c;
assign _c_characterGenerator8x16[567] = 8'h6c;
assign _c_characterGenerator8x16[568] = 8'h6c;
assign _c_characterGenerator8x16[569] = 8'hfe;
assign _c_characterGenerator8x16[570] = 8'h6c;
assign _c_characterGenerator8x16[571] = 8'h6c;
assign _c_characterGenerator8x16[572] = 8'h00;
assign _c_characterGenerator8x16[573] = 8'h00;
assign _c_characterGenerator8x16[574] = 8'h00;
assign _c_characterGenerator8x16[575] = 8'h00;
assign _c_characterGenerator8x16[576] = 8'h18;
assign _c_characterGenerator8x16[577] = 8'h18;
assign _c_characterGenerator8x16[578] = 8'h7c;
assign _c_characterGenerator8x16[579] = 8'hc6;
assign _c_characterGenerator8x16[580] = 8'hc2;
assign _c_characterGenerator8x16[581] = 8'hc0;
assign _c_characterGenerator8x16[582] = 8'h7c;
assign _c_characterGenerator8x16[583] = 8'h06;
assign _c_characterGenerator8x16[584] = 8'h06;
assign _c_characterGenerator8x16[585] = 8'h86;
assign _c_characterGenerator8x16[586] = 8'hc6;
assign _c_characterGenerator8x16[587] = 8'h7c;
assign _c_characterGenerator8x16[588] = 8'h18;
assign _c_characterGenerator8x16[589] = 8'h18;
assign _c_characterGenerator8x16[590] = 8'h00;
assign _c_characterGenerator8x16[591] = 8'h00;
assign _c_characterGenerator8x16[592] = 8'h00;
assign _c_characterGenerator8x16[593] = 8'h00;
assign _c_characterGenerator8x16[594] = 8'h00;
assign _c_characterGenerator8x16[595] = 8'h00;
assign _c_characterGenerator8x16[596] = 8'hc2;
assign _c_characterGenerator8x16[597] = 8'hc6;
assign _c_characterGenerator8x16[598] = 8'h0c;
assign _c_characterGenerator8x16[599] = 8'h18;
assign _c_characterGenerator8x16[600] = 8'h30;
assign _c_characterGenerator8x16[601] = 8'h60;
assign _c_characterGenerator8x16[602] = 8'hc6;
assign _c_characterGenerator8x16[603] = 8'h86;
assign _c_characterGenerator8x16[604] = 8'h00;
assign _c_characterGenerator8x16[605] = 8'h00;
assign _c_characterGenerator8x16[606] = 8'h00;
assign _c_characterGenerator8x16[607] = 8'h00;
assign _c_characterGenerator8x16[608] = 8'h00;
assign _c_characterGenerator8x16[609] = 8'h00;
assign _c_characterGenerator8x16[610] = 8'h38;
assign _c_characterGenerator8x16[611] = 8'h6c;
assign _c_characterGenerator8x16[612] = 8'h6c;
assign _c_characterGenerator8x16[613] = 8'h38;
assign _c_characterGenerator8x16[614] = 8'h76;
assign _c_characterGenerator8x16[615] = 8'hdc;
assign _c_characterGenerator8x16[616] = 8'hcc;
assign _c_characterGenerator8x16[617] = 8'hcc;
assign _c_characterGenerator8x16[618] = 8'hcc;
assign _c_characterGenerator8x16[619] = 8'h76;
assign _c_characterGenerator8x16[620] = 8'h00;
assign _c_characterGenerator8x16[621] = 8'h00;
assign _c_characterGenerator8x16[622] = 8'h00;
assign _c_characterGenerator8x16[623] = 8'h00;
assign _c_characterGenerator8x16[624] = 8'h00;
assign _c_characterGenerator8x16[625] = 8'h30;
assign _c_characterGenerator8x16[626] = 8'h30;
assign _c_characterGenerator8x16[627] = 8'h30;
assign _c_characterGenerator8x16[628] = 8'h60;
assign _c_characterGenerator8x16[629] = 8'h00;
assign _c_characterGenerator8x16[630] = 8'h00;
assign _c_characterGenerator8x16[631] = 8'h00;
assign _c_characterGenerator8x16[632] = 8'h00;
assign _c_characterGenerator8x16[633] = 8'h00;
assign _c_characterGenerator8x16[634] = 8'h00;
assign _c_characterGenerator8x16[635] = 8'h00;
assign _c_characterGenerator8x16[636] = 8'h00;
assign _c_characterGenerator8x16[637] = 8'h00;
assign _c_characterGenerator8x16[638] = 8'h00;
assign _c_characterGenerator8x16[639] = 8'h00;
assign _c_characterGenerator8x16[640] = 8'h00;
assign _c_characterGenerator8x16[641] = 8'h00;
assign _c_characterGenerator8x16[642] = 8'h0c;
assign _c_characterGenerator8x16[643] = 8'h18;
assign _c_characterGenerator8x16[644] = 8'h30;
assign _c_characterGenerator8x16[645] = 8'h30;
assign _c_characterGenerator8x16[646] = 8'h30;
assign _c_characterGenerator8x16[647] = 8'h30;
assign _c_characterGenerator8x16[648] = 8'h30;
assign _c_characterGenerator8x16[649] = 8'h30;
assign _c_characterGenerator8x16[650] = 8'h18;
assign _c_characterGenerator8x16[651] = 8'h0c;
assign _c_characterGenerator8x16[652] = 8'h00;
assign _c_characterGenerator8x16[653] = 8'h00;
assign _c_characterGenerator8x16[654] = 8'h00;
assign _c_characterGenerator8x16[655] = 8'h00;
assign _c_characterGenerator8x16[656] = 8'h00;
assign _c_characterGenerator8x16[657] = 8'h00;
assign _c_characterGenerator8x16[658] = 8'h30;
assign _c_characterGenerator8x16[659] = 8'h18;
assign _c_characterGenerator8x16[660] = 8'h0c;
assign _c_characterGenerator8x16[661] = 8'h0c;
assign _c_characterGenerator8x16[662] = 8'h0c;
assign _c_characterGenerator8x16[663] = 8'h0c;
assign _c_characterGenerator8x16[664] = 8'h0c;
assign _c_characterGenerator8x16[665] = 8'h0c;
assign _c_characterGenerator8x16[666] = 8'h18;
assign _c_characterGenerator8x16[667] = 8'h30;
assign _c_characterGenerator8x16[668] = 8'h00;
assign _c_characterGenerator8x16[669] = 8'h00;
assign _c_characterGenerator8x16[670] = 8'h00;
assign _c_characterGenerator8x16[671] = 8'h00;
assign _c_characterGenerator8x16[672] = 8'h00;
assign _c_characterGenerator8x16[673] = 8'h00;
assign _c_characterGenerator8x16[674] = 8'h00;
assign _c_characterGenerator8x16[675] = 8'h00;
assign _c_characterGenerator8x16[676] = 8'h00;
assign _c_characterGenerator8x16[677] = 8'h66;
assign _c_characterGenerator8x16[678] = 8'h3c;
assign _c_characterGenerator8x16[679] = 8'hff;
assign _c_characterGenerator8x16[680] = 8'h3c;
assign _c_characterGenerator8x16[681] = 8'h66;
assign _c_characterGenerator8x16[682] = 8'h00;
assign _c_characterGenerator8x16[683] = 8'h00;
assign _c_characterGenerator8x16[684] = 8'h00;
assign _c_characterGenerator8x16[685] = 8'h00;
assign _c_characterGenerator8x16[686] = 8'h00;
assign _c_characterGenerator8x16[687] = 8'h00;
assign _c_characterGenerator8x16[688] = 8'h00;
assign _c_characterGenerator8x16[689] = 8'h00;
assign _c_characterGenerator8x16[690] = 8'h00;
assign _c_characterGenerator8x16[691] = 8'h00;
assign _c_characterGenerator8x16[692] = 8'h00;
assign _c_characterGenerator8x16[693] = 8'h18;
assign _c_characterGenerator8x16[694] = 8'h18;
assign _c_characterGenerator8x16[695] = 8'h7e;
assign _c_characterGenerator8x16[696] = 8'h18;
assign _c_characterGenerator8x16[697] = 8'h18;
assign _c_characterGenerator8x16[698] = 8'h00;
assign _c_characterGenerator8x16[699] = 8'h00;
assign _c_characterGenerator8x16[700] = 8'h00;
assign _c_characterGenerator8x16[701] = 8'h00;
assign _c_characterGenerator8x16[702] = 8'h00;
assign _c_characterGenerator8x16[703] = 8'h00;
assign _c_characterGenerator8x16[704] = 8'h00;
assign _c_characterGenerator8x16[705] = 8'h00;
assign _c_characterGenerator8x16[706] = 8'h00;
assign _c_characterGenerator8x16[707] = 8'h00;
assign _c_characterGenerator8x16[708] = 8'h00;
assign _c_characterGenerator8x16[709] = 8'h00;
assign _c_characterGenerator8x16[710] = 8'h00;
assign _c_characterGenerator8x16[711] = 8'h00;
assign _c_characterGenerator8x16[712] = 8'h00;
assign _c_characterGenerator8x16[713] = 8'h18;
assign _c_characterGenerator8x16[714] = 8'h18;
assign _c_characterGenerator8x16[715] = 8'h18;
assign _c_characterGenerator8x16[716] = 8'h30;
assign _c_characterGenerator8x16[717] = 8'h00;
assign _c_characterGenerator8x16[718] = 8'h00;
assign _c_characterGenerator8x16[719] = 8'h00;
assign _c_characterGenerator8x16[720] = 8'h00;
assign _c_characterGenerator8x16[721] = 8'h00;
assign _c_characterGenerator8x16[722] = 8'h00;
assign _c_characterGenerator8x16[723] = 8'h00;
assign _c_characterGenerator8x16[724] = 8'h00;
assign _c_characterGenerator8x16[725] = 8'h00;
assign _c_characterGenerator8x16[726] = 8'h00;
assign _c_characterGenerator8x16[727] = 8'hfe;
assign _c_characterGenerator8x16[728] = 8'h00;
assign _c_characterGenerator8x16[729] = 8'h00;
assign _c_characterGenerator8x16[730] = 8'h00;
assign _c_characterGenerator8x16[731] = 8'h00;
assign _c_characterGenerator8x16[732] = 8'h00;
assign _c_characterGenerator8x16[733] = 8'h00;
assign _c_characterGenerator8x16[734] = 8'h00;
assign _c_characterGenerator8x16[735] = 8'h00;
assign _c_characterGenerator8x16[736] = 8'h00;
assign _c_characterGenerator8x16[737] = 8'h00;
assign _c_characterGenerator8x16[738] = 8'h00;
assign _c_characterGenerator8x16[739] = 8'h00;
assign _c_characterGenerator8x16[740] = 8'h00;
assign _c_characterGenerator8x16[741] = 8'h00;
assign _c_characterGenerator8x16[742] = 8'h00;
assign _c_characterGenerator8x16[743] = 8'h00;
assign _c_characterGenerator8x16[744] = 8'h00;
assign _c_characterGenerator8x16[745] = 8'h00;
assign _c_characterGenerator8x16[746] = 8'h18;
assign _c_characterGenerator8x16[747] = 8'h18;
assign _c_characterGenerator8x16[748] = 8'h00;
assign _c_characterGenerator8x16[749] = 8'h00;
assign _c_characterGenerator8x16[750] = 8'h00;
assign _c_characterGenerator8x16[751] = 8'h00;
assign _c_characterGenerator8x16[752] = 8'h00;
assign _c_characterGenerator8x16[753] = 8'h00;
assign _c_characterGenerator8x16[754] = 8'h00;
assign _c_characterGenerator8x16[755] = 8'h00;
assign _c_characterGenerator8x16[756] = 8'h02;
assign _c_characterGenerator8x16[757] = 8'h06;
assign _c_characterGenerator8x16[758] = 8'h0c;
assign _c_characterGenerator8x16[759] = 8'h18;
assign _c_characterGenerator8x16[760] = 8'h30;
assign _c_characterGenerator8x16[761] = 8'h60;
assign _c_characterGenerator8x16[762] = 8'hc0;
assign _c_characterGenerator8x16[763] = 8'h80;
assign _c_characterGenerator8x16[764] = 8'h00;
assign _c_characterGenerator8x16[765] = 8'h00;
assign _c_characterGenerator8x16[766] = 8'h00;
assign _c_characterGenerator8x16[767] = 8'h00;
assign _c_characterGenerator8x16[768] = 8'h00;
assign _c_characterGenerator8x16[769] = 8'h00;
assign _c_characterGenerator8x16[770] = 8'h38;
assign _c_characterGenerator8x16[771] = 8'h6c;
assign _c_characterGenerator8x16[772] = 8'hc6;
assign _c_characterGenerator8x16[773] = 8'hc6;
assign _c_characterGenerator8x16[774] = 8'hd6;
assign _c_characterGenerator8x16[775] = 8'hd6;
assign _c_characterGenerator8x16[776] = 8'hc6;
assign _c_characterGenerator8x16[777] = 8'hc6;
assign _c_characterGenerator8x16[778] = 8'h6c;
assign _c_characterGenerator8x16[779] = 8'h38;
assign _c_characterGenerator8x16[780] = 8'h00;
assign _c_characterGenerator8x16[781] = 8'h00;
assign _c_characterGenerator8x16[782] = 8'h00;
assign _c_characterGenerator8x16[783] = 8'h00;
assign _c_characterGenerator8x16[784] = 8'h00;
assign _c_characterGenerator8x16[785] = 8'h00;
assign _c_characterGenerator8x16[786] = 8'h18;
assign _c_characterGenerator8x16[787] = 8'h38;
assign _c_characterGenerator8x16[788] = 8'h78;
assign _c_characterGenerator8x16[789] = 8'h18;
assign _c_characterGenerator8x16[790] = 8'h18;
assign _c_characterGenerator8x16[791] = 8'h18;
assign _c_characterGenerator8x16[792] = 8'h18;
assign _c_characterGenerator8x16[793] = 8'h18;
assign _c_characterGenerator8x16[794] = 8'h18;
assign _c_characterGenerator8x16[795] = 8'h7e;
assign _c_characterGenerator8x16[796] = 8'h00;
assign _c_characterGenerator8x16[797] = 8'h00;
assign _c_characterGenerator8x16[798] = 8'h00;
assign _c_characterGenerator8x16[799] = 8'h00;
assign _c_characterGenerator8x16[800] = 8'h00;
assign _c_characterGenerator8x16[801] = 8'h00;
assign _c_characterGenerator8x16[802] = 8'h7c;
assign _c_characterGenerator8x16[803] = 8'hc6;
assign _c_characterGenerator8x16[804] = 8'h06;
assign _c_characterGenerator8x16[805] = 8'h0c;
assign _c_characterGenerator8x16[806] = 8'h18;
assign _c_characterGenerator8x16[807] = 8'h30;
assign _c_characterGenerator8x16[808] = 8'h60;
assign _c_characterGenerator8x16[809] = 8'hc0;
assign _c_characterGenerator8x16[810] = 8'hc6;
assign _c_characterGenerator8x16[811] = 8'hfe;
assign _c_characterGenerator8x16[812] = 8'h00;
assign _c_characterGenerator8x16[813] = 8'h00;
assign _c_characterGenerator8x16[814] = 8'h00;
assign _c_characterGenerator8x16[815] = 8'h00;
assign _c_characterGenerator8x16[816] = 8'h00;
assign _c_characterGenerator8x16[817] = 8'h00;
assign _c_characterGenerator8x16[818] = 8'h7c;
assign _c_characterGenerator8x16[819] = 8'hc6;
assign _c_characterGenerator8x16[820] = 8'h06;
assign _c_characterGenerator8x16[821] = 8'h06;
assign _c_characterGenerator8x16[822] = 8'h3c;
assign _c_characterGenerator8x16[823] = 8'h06;
assign _c_characterGenerator8x16[824] = 8'h06;
assign _c_characterGenerator8x16[825] = 8'h06;
assign _c_characterGenerator8x16[826] = 8'hc6;
assign _c_characterGenerator8x16[827] = 8'h7c;
assign _c_characterGenerator8x16[828] = 8'h00;
assign _c_characterGenerator8x16[829] = 8'h00;
assign _c_characterGenerator8x16[830] = 8'h00;
assign _c_characterGenerator8x16[831] = 8'h00;
assign _c_characterGenerator8x16[832] = 8'h00;
assign _c_characterGenerator8x16[833] = 8'h00;
assign _c_characterGenerator8x16[834] = 8'h0c;
assign _c_characterGenerator8x16[835] = 8'h1c;
assign _c_characterGenerator8x16[836] = 8'h3c;
assign _c_characterGenerator8x16[837] = 8'h6c;
assign _c_characterGenerator8x16[838] = 8'hcc;
assign _c_characterGenerator8x16[839] = 8'hfe;
assign _c_characterGenerator8x16[840] = 8'h0c;
assign _c_characterGenerator8x16[841] = 8'h0c;
assign _c_characterGenerator8x16[842] = 8'h0c;
assign _c_characterGenerator8x16[843] = 8'h1e;
assign _c_characterGenerator8x16[844] = 8'h00;
assign _c_characterGenerator8x16[845] = 8'h00;
assign _c_characterGenerator8x16[846] = 8'h00;
assign _c_characterGenerator8x16[847] = 8'h00;
assign _c_characterGenerator8x16[848] = 8'h00;
assign _c_characterGenerator8x16[849] = 8'h00;
assign _c_characterGenerator8x16[850] = 8'hfe;
assign _c_characterGenerator8x16[851] = 8'hc0;
assign _c_characterGenerator8x16[852] = 8'hc0;
assign _c_characterGenerator8x16[853] = 8'hc0;
assign _c_characterGenerator8x16[854] = 8'hfc;
assign _c_characterGenerator8x16[855] = 8'h06;
assign _c_characterGenerator8x16[856] = 8'h06;
assign _c_characterGenerator8x16[857] = 8'h06;
assign _c_characterGenerator8x16[858] = 8'hc6;
assign _c_characterGenerator8x16[859] = 8'h7c;
assign _c_characterGenerator8x16[860] = 8'h00;
assign _c_characterGenerator8x16[861] = 8'h00;
assign _c_characterGenerator8x16[862] = 8'h00;
assign _c_characterGenerator8x16[863] = 8'h00;
assign _c_characterGenerator8x16[864] = 8'h00;
assign _c_characterGenerator8x16[865] = 8'h00;
assign _c_characterGenerator8x16[866] = 8'h38;
assign _c_characterGenerator8x16[867] = 8'h60;
assign _c_characterGenerator8x16[868] = 8'hc0;
assign _c_characterGenerator8x16[869] = 8'hc0;
assign _c_characterGenerator8x16[870] = 8'hfc;
assign _c_characterGenerator8x16[871] = 8'hc6;
assign _c_characterGenerator8x16[872] = 8'hc6;
assign _c_characterGenerator8x16[873] = 8'hc6;
assign _c_characterGenerator8x16[874] = 8'hc6;
assign _c_characterGenerator8x16[875] = 8'h7c;
assign _c_characterGenerator8x16[876] = 8'h00;
assign _c_characterGenerator8x16[877] = 8'h00;
assign _c_characterGenerator8x16[878] = 8'h00;
assign _c_characterGenerator8x16[879] = 8'h00;
assign _c_characterGenerator8x16[880] = 8'h00;
assign _c_characterGenerator8x16[881] = 8'h00;
assign _c_characterGenerator8x16[882] = 8'hfe;
assign _c_characterGenerator8x16[883] = 8'hc6;
assign _c_characterGenerator8x16[884] = 8'h06;
assign _c_characterGenerator8x16[885] = 8'h06;
assign _c_characterGenerator8x16[886] = 8'h0c;
assign _c_characterGenerator8x16[887] = 8'h18;
assign _c_characterGenerator8x16[888] = 8'h30;
assign _c_characterGenerator8x16[889] = 8'h30;
assign _c_characterGenerator8x16[890] = 8'h30;
assign _c_characterGenerator8x16[891] = 8'h30;
assign _c_characterGenerator8x16[892] = 8'h00;
assign _c_characterGenerator8x16[893] = 8'h00;
assign _c_characterGenerator8x16[894] = 8'h00;
assign _c_characterGenerator8x16[895] = 8'h00;
assign _c_characterGenerator8x16[896] = 8'h00;
assign _c_characterGenerator8x16[897] = 8'h00;
assign _c_characterGenerator8x16[898] = 8'h7c;
assign _c_characterGenerator8x16[899] = 8'hc6;
assign _c_characterGenerator8x16[900] = 8'hc6;
assign _c_characterGenerator8x16[901] = 8'hc6;
assign _c_characterGenerator8x16[902] = 8'h7c;
assign _c_characterGenerator8x16[903] = 8'hc6;
assign _c_characterGenerator8x16[904] = 8'hc6;
assign _c_characterGenerator8x16[905] = 8'hc6;
assign _c_characterGenerator8x16[906] = 8'hc6;
assign _c_characterGenerator8x16[907] = 8'h7c;
assign _c_characterGenerator8x16[908] = 8'h00;
assign _c_characterGenerator8x16[909] = 8'h00;
assign _c_characterGenerator8x16[910] = 8'h00;
assign _c_characterGenerator8x16[911] = 8'h00;
assign _c_characterGenerator8x16[912] = 8'h00;
assign _c_characterGenerator8x16[913] = 8'h00;
assign _c_characterGenerator8x16[914] = 8'h7c;
assign _c_characterGenerator8x16[915] = 8'hc6;
assign _c_characterGenerator8x16[916] = 8'hc6;
assign _c_characterGenerator8x16[917] = 8'hc6;
assign _c_characterGenerator8x16[918] = 8'h7e;
assign _c_characterGenerator8x16[919] = 8'h06;
assign _c_characterGenerator8x16[920] = 8'h06;
assign _c_characterGenerator8x16[921] = 8'h06;
assign _c_characterGenerator8x16[922] = 8'h0c;
assign _c_characterGenerator8x16[923] = 8'h78;
assign _c_characterGenerator8x16[924] = 8'h00;
assign _c_characterGenerator8x16[925] = 8'h00;
assign _c_characterGenerator8x16[926] = 8'h00;
assign _c_characterGenerator8x16[927] = 8'h00;
assign _c_characterGenerator8x16[928] = 8'h00;
assign _c_characterGenerator8x16[929] = 8'h00;
assign _c_characterGenerator8x16[930] = 8'h00;
assign _c_characterGenerator8x16[931] = 8'h00;
assign _c_characterGenerator8x16[932] = 8'h18;
assign _c_characterGenerator8x16[933] = 8'h18;
assign _c_characterGenerator8x16[934] = 8'h00;
assign _c_characterGenerator8x16[935] = 8'h00;
assign _c_characterGenerator8x16[936] = 8'h00;
assign _c_characterGenerator8x16[937] = 8'h18;
assign _c_characterGenerator8x16[938] = 8'h18;
assign _c_characterGenerator8x16[939] = 8'h00;
assign _c_characterGenerator8x16[940] = 8'h00;
assign _c_characterGenerator8x16[941] = 8'h00;
assign _c_characterGenerator8x16[942] = 8'h00;
assign _c_characterGenerator8x16[943] = 8'h00;
assign _c_characterGenerator8x16[944] = 8'h00;
assign _c_characterGenerator8x16[945] = 8'h00;
assign _c_characterGenerator8x16[946] = 8'h00;
assign _c_characterGenerator8x16[947] = 8'h00;
assign _c_characterGenerator8x16[948] = 8'h18;
assign _c_characterGenerator8x16[949] = 8'h18;
assign _c_characterGenerator8x16[950] = 8'h00;
assign _c_characterGenerator8x16[951] = 8'h00;
assign _c_characterGenerator8x16[952] = 8'h00;
assign _c_characterGenerator8x16[953] = 8'h18;
assign _c_characterGenerator8x16[954] = 8'h18;
assign _c_characterGenerator8x16[955] = 8'h30;
assign _c_characterGenerator8x16[956] = 8'h00;
assign _c_characterGenerator8x16[957] = 8'h00;
assign _c_characterGenerator8x16[958] = 8'h00;
assign _c_characterGenerator8x16[959] = 8'h00;
assign _c_characterGenerator8x16[960] = 8'h00;
assign _c_characterGenerator8x16[961] = 8'h00;
assign _c_characterGenerator8x16[962] = 8'h00;
assign _c_characterGenerator8x16[963] = 8'h06;
assign _c_characterGenerator8x16[964] = 8'h0c;
assign _c_characterGenerator8x16[965] = 8'h18;
assign _c_characterGenerator8x16[966] = 8'h30;
assign _c_characterGenerator8x16[967] = 8'h60;
assign _c_characterGenerator8x16[968] = 8'h30;
assign _c_characterGenerator8x16[969] = 8'h18;
assign _c_characterGenerator8x16[970] = 8'h0c;
assign _c_characterGenerator8x16[971] = 8'h06;
assign _c_characterGenerator8x16[972] = 8'h00;
assign _c_characterGenerator8x16[973] = 8'h00;
assign _c_characterGenerator8x16[974] = 8'h00;
assign _c_characterGenerator8x16[975] = 8'h00;
assign _c_characterGenerator8x16[976] = 8'h00;
assign _c_characterGenerator8x16[977] = 8'h00;
assign _c_characterGenerator8x16[978] = 8'h00;
assign _c_characterGenerator8x16[979] = 8'h00;
assign _c_characterGenerator8x16[980] = 8'h00;
assign _c_characterGenerator8x16[981] = 8'h7e;
assign _c_characterGenerator8x16[982] = 8'h00;
assign _c_characterGenerator8x16[983] = 8'h00;
assign _c_characterGenerator8x16[984] = 8'h7e;
assign _c_characterGenerator8x16[985] = 8'h00;
assign _c_characterGenerator8x16[986] = 8'h00;
assign _c_characterGenerator8x16[987] = 8'h00;
assign _c_characterGenerator8x16[988] = 8'h00;
assign _c_characterGenerator8x16[989] = 8'h00;
assign _c_characterGenerator8x16[990] = 8'h00;
assign _c_characterGenerator8x16[991] = 8'h00;
assign _c_characterGenerator8x16[992] = 8'h00;
assign _c_characterGenerator8x16[993] = 8'h00;
assign _c_characterGenerator8x16[994] = 8'h00;
assign _c_characterGenerator8x16[995] = 8'h60;
assign _c_characterGenerator8x16[996] = 8'h30;
assign _c_characterGenerator8x16[997] = 8'h18;
assign _c_characterGenerator8x16[998] = 8'h0c;
assign _c_characterGenerator8x16[999] = 8'h06;
assign _c_characterGenerator8x16[1000] = 8'h0c;
assign _c_characterGenerator8x16[1001] = 8'h18;
assign _c_characterGenerator8x16[1002] = 8'h30;
assign _c_characterGenerator8x16[1003] = 8'h60;
assign _c_characterGenerator8x16[1004] = 8'h00;
assign _c_characterGenerator8x16[1005] = 8'h00;
assign _c_characterGenerator8x16[1006] = 8'h00;
assign _c_characterGenerator8x16[1007] = 8'h00;
assign _c_characterGenerator8x16[1008] = 8'h00;
assign _c_characterGenerator8x16[1009] = 8'h00;
assign _c_characterGenerator8x16[1010] = 8'h7c;
assign _c_characterGenerator8x16[1011] = 8'hc6;
assign _c_characterGenerator8x16[1012] = 8'hc6;
assign _c_characterGenerator8x16[1013] = 8'h0c;
assign _c_characterGenerator8x16[1014] = 8'h18;
assign _c_characterGenerator8x16[1015] = 8'h18;
assign _c_characterGenerator8x16[1016] = 8'h18;
assign _c_characterGenerator8x16[1017] = 8'h00;
assign _c_characterGenerator8x16[1018] = 8'h18;
assign _c_characterGenerator8x16[1019] = 8'h18;
assign _c_characterGenerator8x16[1020] = 8'h00;
assign _c_characterGenerator8x16[1021] = 8'h00;
assign _c_characterGenerator8x16[1022] = 8'h00;
assign _c_characterGenerator8x16[1023] = 8'h00;
assign _c_characterGenerator8x16[1024] = 8'h00;
assign _c_characterGenerator8x16[1025] = 8'h00;
assign _c_characterGenerator8x16[1026] = 8'h00;
assign _c_characterGenerator8x16[1027] = 8'h7c;
assign _c_characterGenerator8x16[1028] = 8'hc6;
assign _c_characterGenerator8x16[1029] = 8'hc6;
assign _c_characterGenerator8x16[1030] = 8'hde;
assign _c_characterGenerator8x16[1031] = 8'hde;
assign _c_characterGenerator8x16[1032] = 8'hde;
assign _c_characterGenerator8x16[1033] = 8'hdc;
assign _c_characterGenerator8x16[1034] = 8'hc0;
assign _c_characterGenerator8x16[1035] = 8'h7c;
assign _c_characterGenerator8x16[1036] = 8'h00;
assign _c_characterGenerator8x16[1037] = 8'h00;
assign _c_characterGenerator8x16[1038] = 8'h00;
assign _c_characterGenerator8x16[1039] = 8'h00;
assign _c_characterGenerator8x16[1040] = 8'h00;
assign _c_characterGenerator8x16[1041] = 8'h00;
assign _c_characterGenerator8x16[1042] = 8'h10;
assign _c_characterGenerator8x16[1043] = 8'h38;
assign _c_characterGenerator8x16[1044] = 8'h6c;
assign _c_characterGenerator8x16[1045] = 8'hc6;
assign _c_characterGenerator8x16[1046] = 8'hc6;
assign _c_characterGenerator8x16[1047] = 8'hfe;
assign _c_characterGenerator8x16[1048] = 8'hc6;
assign _c_characterGenerator8x16[1049] = 8'hc6;
assign _c_characterGenerator8x16[1050] = 8'hc6;
assign _c_characterGenerator8x16[1051] = 8'hc6;
assign _c_characterGenerator8x16[1052] = 8'h00;
assign _c_characterGenerator8x16[1053] = 8'h00;
assign _c_characterGenerator8x16[1054] = 8'h00;
assign _c_characterGenerator8x16[1055] = 8'h00;
assign _c_characterGenerator8x16[1056] = 8'h00;
assign _c_characterGenerator8x16[1057] = 8'h00;
assign _c_characterGenerator8x16[1058] = 8'hfc;
assign _c_characterGenerator8x16[1059] = 8'h66;
assign _c_characterGenerator8x16[1060] = 8'h66;
assign _c_characterGenerator8x16[1061] = 8'h66;
assign _c_characterGenerator8x16[1062] = 8'h7c;
assign _c_characterGenerator8x16[1063] = 8'h66;
assign _c_characterGenerator8x16[1064] = 8'h66;
assign _c_characterGenerator8x16[1065] = 8'h66;
assign _c_characterGenerator8x16[1066] = 8'h66;
assign _c_characterGenerator8x16[1067] = 8'hfc;
assign _c_characterGenerator8x16[1068] = 8'h00;
assign _c_characterGenerator8x16[1069] = 8'h00;
assign _c_characterGenerator8x16[1070] = 8'h00;
assign _c_characterGenerator8x16[1071] = 8'h00;
assign _c_characterGenerator8x16[1072] = 8'h00;
assign _c_characterGenerator8x16[1073] = 8'h00;
assign _c_characterGenerator8x16[1074] = 8'h3c;
assign _c_characterGenerator8x16[1075] = 8'h66;
assign _c_characterGenerator8x16[1076] = 8'hc2;
assign _c_characterGenerator8x16[1077] = 8'hc0;
assign _c_characterGenerator8x16[1078] = 8'hc0;
assign _c_characterGenerator8x16[1079] = 8'hc0;
assign _c_characterGenerator8x16[1080] = 8'hc0;
assign _c_characterGenerator8x16[1081] = 8'hc2;
assign _c_characterGenerator8x16[1082] = 8'h66;
assign _c_characterGenerator8x16[1083] = 8'h3c;
assign _c_characterGenerator8x16[1084] = 8'h00;
assign _c_characterGenerator8x16[1085] = 8'h00;
assign _c_characterGenerator8x16[1086] = 8'h00;
assign _c_characterGenerator8x16[1087] = 8'h00;
assign _c_characterGenerator8x16[1088] = 8'h00;
assign _c_characterGenerator8x16[1089] = 8'h00;
assign _c_characterGenerator8x16[1090] = 8'hf8;
assign _c_characterGenerator8x16[1091] = 8'h6c;
assign _c_characterGenerator8x16[1092] = 8'h66;
assign _c_characterGenerator8x16[1093] = 8'h66;
assign _c_characterGenerator8x16[1094] = 8'h66;
assign _c_characterGenerator8x16[1095] = 8'h66;
assign _c_characterGenerator8x16[1096] = 8'h66;
assign _c_characterGenerator8x16[1097] = 8'h66;
assign _c_characterGenerator8x16[1098] = 8'h6c;
assign _c_characterGenerator8x16[1099] = 8'hf8;
assign _c_characterGenerator8x16[1100] = 8'h00;
assign _c_characterGenerator8x16[1101] = 8'h00;
assign _c_characterGenerator8x16[1102] = 8'h00;
assign _c_characterGenerator8x16[1103] = 8'h00;
assign _c_characterGenerator8x16[1104] = 8'h00;
assign _c_characterGenerator8x16[1105] = 8'h00;
assign _c_characterGenerator8x16[1106] = 8'hfe;
assign _c_characterGenerator8x16[1107] = 8'h66;
assign _c_characterGenerator8x16[1108] = 8'h62;
assign _c_characterGenerator8x16[1109] = 8'h68;
assign _c_characterGenerator8x16[1110] = 8'h78;
assign _c_characterGenerator8x16[1111] = 8'h68;
assign _c_characterGenerator8x16[1112] = 8'h60;
assign _c_characterGenerator8x16[1113] = 8'h62;
assign _c_characterGenerator8x16[1114] = 8'h66;
assign _c_characterGenerator8x16[1115] = 8'hfe;
assign _c_characterGenerator8x16[1116] = 8'h00;
assign _c_characterGenerator8x16[1117] = 8'h00;
assign _c_characterGenerator8x16[1118] = 8'h00;
assign _c_characterGenerator8x16[1119] = 8'h00;
assign _c_characterGenerator8x16[1120] = 8'h00;
assign _c_characterGenerator8x16[1121] = 8'h00;
assign _c_characterGenerator8x16[1122] = 8'hfe;
assign _c_characterGenerator8x16[1123] = 8'h66;
assign _c_characterGenerator8x16[1124] = 8'h62;
assign _c_characterGenerator8x16[1125] = 8'h68;
assign _c_characterGenerator8x16[1126] = 8'h78;
assign _c_characterGenerator8x16[1127] = 8'h68;
assign _c_characterGenerator8x16[1128] = 8'h60;
assign _c_characterGenerator8x16[1129] = 8'h60;
assign _c_characterGenerator8x16[1130] = 8'h60;
assign _c_characterGenerator8x16[1131] = 8'hf0;
assign _c_characterGenerator8x16[1132] = 8'h00;
assign _c_characterGenerator8x16[1133] = 8'h00;
assign _c_characterGenerator8x16[1134] = 8'h00;
assign _c_characterGenerator8x16[1135] = 8'h00;
assign _c_characterGenerator8x16[1136] = 8'h00;
assign _c_characterGenerator8x16[1137] = 8'h00;
assign _c_characterGenerator8x16[1138] = 8'h3c;
assign _c_characterGenerator8x16[1139] = 8'h66;
assign _c_characterGenerator8x16[1140] = 8'hc2;
assign _c_characterGenerator8x16[1141] = 8'hc0;
assign _c_characterGenerator8x16[1142] = 8'hc0;
assign _c_characterGenerator8x16[1143] = 8'hde;
assign _c_characterGenerator8x16[1144] = 8'hc6;
assign _c_characterGenerator8x16[1145] = 8'hc6;
assign _c_characterGenerator8x16[1146] = 8'h66;
assign _c_characterGenerator8x16[1147] = 8'h3a;
assign _c_characterGenerator8x16[1148] = 8'h00;
assign _c_characterGenerator8x16[1149] = 8'h00;
assign _c_characterGenerator8x16[1150] = 8'h00;
assign _c_characterGenerator8x16[1151] = 8'h00;
assign _c_characterGenerator8x16[1152] = 8'h00;
assign _c_characterGenerator8x16[1153] = 8'h00;
assign _c_characterGenerator8x16[1154] = 8'hc6;
assign _c_characterGenerator8x16[1155] = 8'hc6;
assign _c_characterGenerator8x16[1156] = 8'hc6;
assign _c_characterGenerator8x16[1157] = 8'hc6;
assign _c_characterGenerator8x16[1158] = 8'hfe;
assign _c_characterGenerator8x16[1159] = 8'hc6;
assign _c_characterGenerator8x16[1160] = 8'hc6;
assign _c_characterGenerator8x16[1161] = 8'hc6;
assign _c_characterGenerator8x16[1162] = 8'hc6;
assign _c_characterGenerator8x16[1163] = 8'hc6;
assign _c_characterGenerator8x16[1164] = 8'h00;
assign _c_characterGenerator8x16[1165] = 8'h00;
assign _c_characterGenerator8x16[1166] = 8'h00;
assign _c_characterGenerator8x16[1167] = 8'h00;
assign _c_characterGenerator8x16[1168] = 8'h00;
assign _c_characterGenerator8x16[1169] = 8'h00;
assign _c_characterGenerator8x16[1170] = 8'h3c;
assign _c_characterGenerator8x16[1171] = 8'h18;
assign _c_characterGenerator8x16[1172] = 8'h18;
assign _c_characterGenerator8x16[1173] = 8'h18;
assign _c_characterGenerator8x16[1174] = 8'h18;
assign _c_characterGenerator8x16[1175] = 8'h18;
assign _c_characterGenerator8x16[1176] = 8'h18;
assign _c_characterGenerator8x16[1177] = 8'h18;
assign _c_characterGenerator8x16[1178] = 8'h18;
assign _c_characterGenerator8x16[1179] = 8'h3c;
assign _c_characterGenerator8x16[1180] = 8'h00;
assign _c_characterGenerator8x16[1181] = 8'h00;
assign _c_characterGenerator8x16[1182] = 8'h00;
assign _c_characterGenerator8x16[1183] = 8'h00;
assign _c_characterGenerator8x16[1184] = 8'h00;
assign _c_characterGenerator8x16[1185] = 8'h00;
assign _c_characterGenerator8x16[1186] = 8'h1e;
assign _c_characterGenerator8x16[1187] = 8'h0c;
assign _c_characterGenerator8x16[1188] = 8'h0c;
assign _c_characterGenerator8x16[1189] = 8'h0c;
assign _c_characterGenerator8x16[1190] = 8'h0c;
assign _c_characterGenerator8x16[1191] = 8'h0c;
assign _c_characterGenerator8x16[1192] = 8'hcc;
assign _c_characterGenerator8x16[1193] = 8'hcc;
assign _c_characterGenerator8x16[1194] = 8'hcc;
assign _c_characterGenerator8x16[1195] = 8'h78;
assign _c_characterGenerator8x16[1196] = 8'h00;
assign _c_characterGenerator8x16[1197] = 8'h00;
assign _c_characterGenerator8x16[1198] = 8'h00;
assign _c_characterGenerator8x16[1199] = 8'h00;
assign _c_characterGenerator8x16[1200] = 8'h00;
assign _c_characterGenerator8x16[1201] = 8'h00;
assign _c_characterGenerator8x16[1202] = 8'he6;
assign _c_characterGenerator8x16[1203] = 8'h66;
assign _c_characterGenerator8x16[1204] = 8'h66;
assign _c_characterGenerator8x16[1205] = 8'h6c;
assign _c_characterGenerator8x16[1206] = 8'h78;
assign _c_characterGenerator8x16[1207] = 8'h78;
assign _c_characterGenerator8x16[1208] = 8'h6c;
assign _c_characterGenerator8x16[1209] = 8'h66;
assign _c_characterGenerator8x16[1210] = 8'h66;
assign _c_characterGenerator8x16[1211] = 8'he6;
assign _c_characterGenerator8x16[1212] = 8'h00;
assign _c_characterGenerator8x16[1213] = 8'h00;
assign _c_characterGenerator8x16[1214] = 8'h00;
assign _c_characterGenerator8x16[1215] = 8'h00;
assign _c_characterGenerator8x16[1216] = 8'h00;
assign _c_characterGenerator8x16[1217] = 8'h00;
assign _c_characterGenerator8x16[1218] = 8'hf0;
assign _c_characterGenerator8x16[1219] = 8'h60;
assign _c_characterGenerator8x16[1220] = 8'h60;
assign _c_characterGenerator8x16[1221] = 8'h60;
assign _c_characterGenerator8x16[1222] = 8'h60;
assign _c_characterGenerator8x16[1223] = 8'h60;
assign _c_characterGenerator8x16[1224] = 8'h60;
assign _c_characterGenerator8x16[1225] = 8'h62;
assign _c_characterGenerator8x16[1226] = 8'h66;
assign _c_characterGenerator8x16[1227] = 8'hfe;
assign _c_characterGenerator8x16[1228] = 8'h00;
assign _c_characterGenerator8x16[1229] = 8'h00;
assign _c_characterGenerator8x16[1230] = 8'h00;
assign _c_characterGenerator8x16[1231] = 8'h00;
assign _c_characterGenerator8x16[1232] = 8'h00;
assign _c_characterGenerator8x16[1233] = 8'h00;
assign _c_characterGenerator8x16[1234] = 8'hc6;
assign _c_characterGenerator8x16[1235] = 8'hee;
assign _c_characterGenerator8x16[1236] = 8'hfe;
assign _c_characterGenerator8x16[1237] = 8'hfe;
assign _c_characterGenerator8x16[1238] = 8'hd6;
assign _c_characterGenerator8x16[1239] = 8'hc6;
assign _c_characterGenerator8x16[1240] = 8'hc6;
assign _c_characterGenerator8x16[1241] = 8'hc6;
assign _c_characterGenerator8x16[1242] = 8'hc6;
assign _c_characterGenerator8x16[1243] = 8'hc6;
assign _c_characterGenerator8x16[1244] = 8'h00;
assign _c_characterGenerator8x16[1245] = 8'h00;
assign _c_characterGenerator8x16[1246] = 8'h00;
assign _c_characterGenerator8x16[1247] = 8'h00;
assign _c_characterGenerator8x16[1248] = 8'h00;
assign _c_characterGenerator8x16[1249] = 8'h00;
assign _c_characterGenerator8x16[1250] = 8'hc6;
assign _c_characterGenerator8x16[1251] = 8'he6;
assign _c_characterGenerator8x16[1252] = 8'hf6;
assign _c_characterGenerator8x16[1253] = 8'hfe;
assign _c_characterGenerator8x16[1254] = 8'hde;
assign _c_characterGenerator8x16[1255] = 8'hce;
assign _c_characterGenerator8x16[1256] = 8'hc6;
assign _c_characterGenerator8x16[1257] = 8'hc6;
assign _c_characterGenerator8x16[1258] = 8'hc6;
assign _c_characterGenerator8x16[1259] = 8'hc6;
assign _c_characterGenerator8x16[1260] = 8'h00;
assign _c_characterGenerator8x16[1261] = 8'h00;
assign _c_characterGenerator8x16[1262] = 8'h00;
assign _c_characterGenerator8x16[1263] = 8'h00;
assign _c_characterGenerator8x16[1264] = 8'h00;
assign _c_characterGenerator8x16[1265] = 8'h00;
assign _c_characterGenerator8x16[1266] = 8'h7c;
assign _c_characterGenerator8x16[1267] = 8'hc6;
assign _c_characterGenerator8x16[1268] = 8'hc6;
assign _c_characterGenerator8x16[1269] = 8'hc6;
assign _c_characterGenerator8x16[1270] = 8'hc6;
assign _c_characterGenerator8x16[1271] = 8'hc6;
assign _c_characterGenerator8x16[1272] = 8'hc6;
assign _c_characterGenerator8x16[1273] = 8'hc6;
assign _c_characterGenerator8x16[1274] = 8'hc6;
assign _c_characterGenerator8x16[1275] = 8'h7c;
assign _c_characterGenerator8x16[1276] = 8'h00;
assign _c_characterGenerator8x16[1277] = 8'h00;
assign _c_characterGenerator8x16[1278] = 8'h00;
assign _c_characterGenerator8x16[1279] = 8'h00;
assign _c_characterGenerator8x16[1280] = 8'h00;
assign _c_characterGenerator8x16[1281] = 8'h00;
assign _c_characterGenerator8x16[1282] = 8'hfc;
assign _c_characterGenerator8x16[1283] = 8'h66;
assign _c_characterGenerator8x16[1284] = 8'h66;
assign _c_characterGenerator8x16[1285] = 8'h66;
assign _c_characterGenerator8x16[1286] = 8'h7c;
assign _c_characterGenerator8x16[1287] = 8'h60;
assign _c_characterGenerator8x16[1288] = 8'h60;
assign _c_characterGenerator8x16[1289] = 8'h60;
assign _c_characterGenerator8x16[1290] = 8'h60;
assign _c_characterGenerator8x16[1291] = 8'hf0;
assign _c_characterGenerator8x16[1292] = 8'h00;
assign _c_characterGenerator8x16[1293] = 8'h00;
assign _c_characterGenerator8x16[1294] = 8'h00;
assign _c_characterGenerator8x16[1295] = 8'h00;
assign _c_characterGenerator8x16[1296] = 8'h00;
assign _c_characterGenerator8x16[1297] = 8'h00;
assign _c_characterGenerator8x16[1298] = 8'h7c;
assign _c_characterGenerator8x16[1299] = 8'hc6;
assign _c_characterGenerator8x16[1300] = 8'hc6;
assign _c_characterGenerator8x16[1301] = 8'hc6;
assign _c_characterGenerator8x16[1302] = 8'hc6;
assign _c_characterGenerator8x16[1303] = 8'hc6;
assign _c_characterGenerator8x16[1304] = 8'hc6;
assign _c_characterGenerator8x16[1305] = 8'hd6;
assign _c_characterGenerator8x16[1306] = 8'hde;
assign _c_characterGenerator8x16[1307] = 8'h7c;
assign _c_characterGenerator8x16[1308] = 8'h0c;
assign _c_characterGenerator8x16[1309] = 8'h0e;
assign _c_characterGenerator8x16[1310] = 8'h00;
assign _c_characterGenerator8x16[1311] = 8'h00;
assign _c_characterGenerator8x16[1312] = 8'h00;
assign _c_characterGenerator8x16[1313] = 8'h00;
assign _c_characterGenerator8x16[1314] = 8'hfc;
assign _c_characterGenerator8x16[1315] = 8'h66;
assign _c_characterGenerator8x16[1316] = 8'h66;
assign _c_characterGenerator8x16[1317] = 8'h66;
assign _c_characterGenerator8x16[1318] = 8'h7c;
assign _c_characterGenerator8x16[1319] = 8'h6c;
assign _c_characterGenerator8x16[1320] = 8'h66;
assign _c_characterGenerator8x16[1321] = 8'h66;
assign _c_characterGenerator8x16[1322] = 8'h66;
assign _c_characterGenerator8x16[1323] = 8'he6;
assign _c_characterGenerator8x16[1324] = 8'h00;
assign _c_characterGenerator8x16[1325] = 8'h00;
assign _c_characterGenerator8x16[1326] = 8'h00;
assign _c_characterGenerator8x16[1327] = 8'h00;
assign _c_characterGenerator8x16[1328] = 8'h00;
assign _c_characterGenerator8x16[1329] = 8'h00;
assign _c_characterGenerator8x16[1330] = 8'h7c;
assign _c_characterGenerator8x16[1331] = 8'hc6;
assign _c_characterGenerator8x16[1332] = 8'hc6;
assign _c_characterGenerator8x16[1333] = 8'h60;
assign _c_characterGenerator8x16[1334] = 8'h38;
assign _c_characterGenerator8x16[1335] = 8'h0c;
assign _c_characterGenerator8x16[1336] = 8'h06;
assign _c_characterGenerator8x16[1337] = 8'hc6;
assign _c_characterGenerator8x16[1338] = 8'hc6;
assign _c_characterGenerator8x16[1339] = 8'h7c;
assign _c_characterGenerator8x16[1340] = 8'h00;
assign _c_characterGenerator8x16[1341] = 8'h00;
assign _c_characterGenerator8x16[1342] = 8'h00;
assign _c_characterGenerator8x16[1343] = 8'h00;
assign _c_characterGenerator8x16[1344] = 8'h00;
assign _c_characterGenerator8x16[1345] = 8'h00;
assign _c_characterGenerator8x16[1346] = 8'h7e;
assign _c_characterGenerator8x16[1347] = 8'h7e;
assign _c_characterGenerator8x16[1348] = 8'h5a;
assign _c_characterGenerator8x16[1349] = 8'h18;
assign _c_characterGenerator8x16[1350] = 8'h18;
assign _c_characterGenerator8x16[1351] = 8'h18;
assign _c_characterGenerator8x16[1352] = 8'h18;
assign _c_characterGenerator8x16[1353] = 8'h18;
assign _c_characterGenerator8x16[1354] = 8'h18;
assign _c_characterGenerator8x16[1355] = 8'h3c;
assign _c_characterGenerator8x16[1356] = 8'h00;
assign _c_characterGenerator8x16[1357] = 8'h00;
assign _c_characterGenerator8x16[1358] = 8'h00;
assign _c_characterGenerator8x16[1359] = 8'h00;
assign _c_characterGenerator8x16[1360] = 8'h00;
assign _c_characterGenerator8x16[1361] = 8'h00;
assign _c_characterGenerator8x16[1362] = 8'hc6;
assign _c_characterGenerator8x16[1363] = 8'hc6;
assign _c_characterGenerator8x16[1364] = 8'hc6;
assign _c_characterGenerator8x16[1365] = 8'hc6;
assign _c_characterGenerator8x16[1366] = 8'hc6;
assign _c_characterGenerator8x16[1367] = 8'hc6;
assign _c_characterGenerator8x16[1368] = 8'hc6;
assign _c_characterGenerator8x16[1369] = 8'hc6;
assign _c_characterGenerator8x16[1370] = 8'hc6;
assign _c_characterGenerator8x16[1371] = 8'h7c;
assign _c_characterGenerator8x16[1372] = 8'h00;
assign _c_characterGenerator8x16[1373] = 8'h00;
assign _c_characterGenerator8x16[1374] = 8'h00;
assign _c_characterGenerator8x16[1375] = 8'h00;
assign _c_characterGenerator8x16[1376] = 8'h00;
assign _c_characterGenerator8x16[1377] = 8'h00;
assign _c_characterGenerator8x16[1378] = 8'hc6;
assign _c_characterGenerator8x16[1379] = 8'hc6;
assign _c_characterGenerator8x16[1380] = 8'hc6;
assign _c_characterGenerator8x16[1381] = 8'hc6;
assign _c_characterGenerator8x16[1382] = 8'hc6;
assign _c_characterGenerator8x16[1383] = 8'hc6;
assign _c_characterGenerator8x16[1384] = 8'hc6;
assign _c_characterGenerator8x16[1385] = 8'h6c;
assign _c_characterGenerator8x16[1386] = 8'h38;
assign _c_characterGenerator8x16[1387] = 8'h10;
assign _c_characterGenerator8x16[1388] = 8'h00;
assign _c_characterGenerator8x16[1389] = 8'h00;
assign _c_characterGenerator8x16[1390] = 8'h00;
assign _c_characterGenerator8x16[1391] = 8'h00;
assign _c_characterGenerator8x16[1392] = 8'h00;
assign _c_characterGenerator8x16[1393] = 8'h00;
assign _c_characterGenerator8x16[1394] = 8'hc6;
assign _c_characterGenerator8x16[1395] = 8'hc6;
assign _c_characterGenerator8x16[1396] = 8'hc6;
assign _c_characterGenerator8x16[1397] = 8'hc6;
assign _c_characterGenerator8x16[1398] = 8'hd6;
assign _c_characterGenerator8x16[1399] = 8'hd6;
assign _c_characterGenerator8x16[1400] = 8'hd6;
assign _c_characterGenerator8x16[1401] = 8'hfe;
assign _c_characterGenerator8x16[1402] = 8'hee;
assign _c_characterGenerator8x16[1403] = 8'h6c;
assign _c_characterGenerator8x16[1404] = 8'h00;
assign _c_characterGenerator8x16[1405] = 8'h00;
assign _c_characterGenerator8x16[1406] = 8'h00;
assign _c_characterGenerator8x16[1407] = 8'h00;
assign _c_characterGenerator8x16[1408] = 8'h00;
assign _c_characterGenerator8x16[1409] = 8'h00;
assign _c_characterGenerator8x16[1410] = 8'hc6;
assign _c_characterGenerator8x16[1411] = 8'hc6;
assign _c_characterGenerator8x16[1412] = 8'h6c;
assign _c_characterGenerator8x16[1413] = 8'h7c;
assign _c_characterGenerator8x16[1414] = 8'h38;
assign _c_characterGenerator8x16[1415] = 8'h38;
assign _c_characterGenerator8x16[1416] = 8'h7c;
assign _c_characterGenerator8x16[1417] = 8'h6c;
assign _c_characterGenerator8x16[1418] = 8'hc6;
assign _c_characterGenerator8x16[1419] = 8'hc6;
assign _c_characterGenerator8x16[1420] = 8'h00;
assign _c_characterGenerator8x16[1421] = 8'h00;
assign _c_characterGenerator8x16[1422] = 8'h00;
assign _c_characterGenerator8x16[1423] = 8'h00;
assign _c_characterGenerator8x16[1424] = 8'h00;
assign _c_characterGenerator8x16[1425] = 8'h00;
assign _c_characterGenerator8x16[1426] = 8'h66;
assign _c_characterGenerator8x16[1427] = 8'h66;
assign _c_characterGenerator8x16[1428] = 8'h66;
assign _c_characterGenerator8x16[1429] = 8'h66;
assign _c_characterGenerator8x16[1430] = 8'h3c;
assign _c_characterGenerator8x16[1431] = 8'h18;
assign _c_characterGenerator8x16[1432] = 8'h18;
assign _c_characterGenerator8x16[1433] = 8'h18;
assign _c_characterGenerator8x16[1434] = 8'h18;
assign _c_characterGenerator8x16[1435] = 8'h3c;
assign _c_characterGenerator8x16[1436] = 8'h00;
assign _c_characterGenerator8x16[1437] = 8'h00;
assign _c_characterGenerator8x16[1438] = 8'h00;
assign _c_characterGenerator8x16[1439] = 8'h00;
assign _c_characterGenerator8x16[1440] = 8'h00;
assign _c_characterGenerator8x16[1441] = 8'h00;
assign _c_characterGenerator8x16[1442] = 8'hfe;
assign _c_characterGenerator8x16[1443] = 8'hc6;
assign _c_characterGenerator8x16[1444] = 8'h86;
assign _c_characterGenerator8x16[1445] = 8'h0c;
assign _c_characterGenerator8x16[1446] = 8'h18;
assign _c_characterGenerator8x16[1447] = 8'h30;
assign _c_characterGenerator8x16[1448] = 8'h60;
assign _c_characterGenerator8x16[1449] = 8'hc2;
assign _c_characterGenerator8x16[1450] = 8'hc6;
assign _c_characterGenerator8x16[1451] = 8'hfe;
assign _c_characterGenerator8x16[1452] = 8'h00;
assign _c_characterGenerator8x16[1453] = 8'h00;
assign _c_characterGenerator8x16[1454] = 8'h00;
assign _c_characterGenerator8x16[1455] = 8'h00;
assign _c_characterGenerator8x16[1456] = 8'h00;
assign _c_characterGenerator8x16[1457] = 8'h00;
assign _c_characterGenerator8x16[1458] = 8'h3c;
assign _c_characterGenerator8x16[1459] = 8'h30;
assign _c_characterGenerator8x16[1460] = 8'h30;
assign _c_characterGenerator8x16[1461] = 8'h30;
assign _c_characterGenerator8x16[1462] = 8'h30;
assign _c_characterGenerator8x16[1463] = 8'h30;
assign _c_characterGenerator8x16[1464] = 8'h30;
assign _c_characterGenerator8x16[1465] = 8'h30;
assign _c_characterGenerator8x16[1466] = 8'h30;
assign _c_characterGenerator8x16[1467] = 8'h3c;
assign _c_characterGenerator8x16[1468] = 8'h00;
assign _c_characterGenerator8x16[1469] = 8'h00;
assign _c_characterGenerator8x16[1470] = 8'h00;
assign _c_characterGenerator8x16[1471] = 8'h00;
assign _c_characterGenerator8x16[1472] = 8'h00;
assign _c_characterGenerator8x16[1473] = 8'h00;
assign _c_characterGenerator8x16[1474] = 8'h00;
assign _c_characterGenerator8x16[1475] = 8'h80;
assign _c_characterGenerator8x16[1476] = 8'hc0;
assign _c_characterGenerator8x16[1477] = 8'he0;
assign _c_characterGenerator8x16[1478] = 8'h70;
assign _c_characterGenerator8x16[1479] = 8'h38;
assign _c_characterGenerator8x16[1480] = 8'h1c;
assign _c_characterGenerator8x16[1481] = 8'h0e;
assign _c_characterGenerator8x16[1482] = 8'h06;
assign _c_characterGenerator8x16[1483] = 8'h02;
assign _c_characterGenerator8x16[1484] = 8'h00;
assign _c_characterGenerator8x16[1485] = 8'h00;
assign _c_characterGenerator8x16[1486] = 8'h00;
assign _c_characterGenerator8x16[1487] = 8'h00;
assign _c_characterGenerator8x16[1488] = 8'h00;
assign _c_characterGenerator8x16[1489] = 8'h00;
assign _c_characterGenerator8x16[1490] = 8'h3c;
assign _c_characterGenerator8x16[1491] = 8'h0c;
assign _c_characterGenerator8x16[1492] = 8'h0c;
assign _c_characterGenerator8x16[1493] = 8'h0c;
assign _c_characterGenerator8x16[1494] = 8'h0c;
assign _c_characterGenerator8x16[1495] = 8'h0c;
assign _c_characterGenerator8x16[1496] = 8'h0c;
assign _c_characterGenerator8x16[1497] = 8'h0c;
assign _c_characterGenerator8x16[1498] = 8'h0c;
assign _c_characterGenerator8x16[1499] = 8'h3c;
assign _c_characterGenerator8x16[1500] = 8'h00;
assign _c_characterGenerator8x16[1501] = 8'h00;
assign _c_characterGenerator8x16[1502] = 8'h00;
assign _c_characterGenerator8x16[1503] = 8'h00;
assign _c_characterGenerator8x16[1504] = 8'h10;
assign _c_characterGenerator8x16[1505] = 8'h38;
assign _c_characterGenerator8x16[1506] = 8'h6c;
assign _c_characterGenerator8x16[1507] = 8'hc6;
assign _c_characterGenerator8x16[1508] = 8'h00;
assign _c_characterGenerator8x16[1509] = 8'h00;
assign _c_characterGenerator8x16[1510] = 8'h00;
assign _c_characterGenerator8x16[1511] = 8'h00;
assign _c_characterGenerator8x16[1512] = 8'h00;
assign _c_characterGenerator8x16[1513] = 8'h00;
assign _c_characterGenerator8x16[1514] = 8'h00;
assign _c_characterGenerator8x16[1515] = 8'h00;
assign _c_characterGenerator8x16[1516] = 8'h00;
assign _c_characterGenerator8x16[1517] = 8'h00;
assign _c_characterGenerator8x16[1518] = 8'h00;
assign _c_characterGenerator8x16[1519] = 8'h00;
assign _c_characterGenerator8x16[1520] = 8'h00;
assign _c_characterGenerator8x16[1521] = 8'h00;
assign _c_characterGenerator8x16[1522] = 8'h00;
assign _c_characterGenerator8x16[1523] = 8'h00;
assign _c_characterGenerator8x16[1524] = 8'h00;
assign _c_characterGenerator8x16[1525] = 8'h00;
assign _c_characterGenerator8x16[1526] = 8'h00;
assign _c_characterGenerator8x16[1527] = 8'h00;
assign _c_characterGenerator8x16[1528] = 8'h00;
assign _c_characterGenerator8x16[1529] = 8'h00;
assign _c_characterGenerator8x16[1530] = 8'h00;
assign _c_characterGenerator8x16[1531] = 8'h00;
assign _c_characterGenerator8x16[1532] = 8'h00;
assign _c_characterGenerator8x16[1533] = 8'hff;
assign _c_characterGenerator8x16[1534] = 8'h00;
assign _c_characterGenerator8x16[1535] = 8'h00;
assign _c_characterGenerator8x16[1536] = 8'h30;
assign _c_characterGenerator8x16[1537] = 8'h30;
assign _c_characterGenerator8x16[1538] = 8'h18;
assign _c_characterGenerator8x16[1539] = 8'h00;
assign _c_characterGenerator8x16[1540] = 8'h00;
assign _c_characterGenerator8x16[1541] = 8'h00;
assign _c_characterGenerator8x16[1542] = 8'h00;
assign _c_characterGenerator8x16[1543] = 8'h00;
assign _c_characterGenerator8x16[1544] = 8'h00;
assign _c_characterGenerator8x16[1545] = 8'h00;
assign _c_characterGenerator8x16[1546] = 8'h00;
assign _c_characterGenerator8x16[1547] = 8'h00;
assign _c_characterGenerator8x16[1548] = 8'h00;
assign _c_characterGenerator8x16[1549] = 8'h00;
assign _c_characterGenerator8x16[1550] = 8'h00;
assign _c_characterGenerator8x16[1551] = 8'h00;
assign _c_characterGenerator8x16[1552] = 8'h00;
assign _c_characterGenerator8x16[1553] = 8'h00;
assign _c_characterGenerator8x16[1554] = 8'h00;
assign _c_characterGenerator8x16[1555] = 8'h00;
assign _c_characterGenerator8x16[1556] = 8'h00;
assign _c_characterGenerator8x16[1557] = 8'h78;
assign _c_characterGenerator8x16[1558] = 8'h0c;
assign _c_characterGenerator8x16[1559] = 8'h7c;
assign _c_characterGenerator8x16[1560] = 8'hcc;
assign _c_characterGenerator8x16[1561] = 8'hcc;
assign _c_characterGenerator8x16[1562] = 8'hcc;
assign _c_characterGenerator8x16[1563] = 8'h76;
assign _c_characterGenerator8x16[1564] = 8'h00;
assign _c_characterGenerator8x16[1565] = 8'h00;
assign _c_characterGenerator8x16[1566] = 8'h00;
assign _c_characterGenerator8x16[1567] = 8'h00;
assign _c_characterGenerator8x16[1568] = 8'h00;
assign _c_characterGenerator8x16[1569] = 8'h00;
assign _c_characterGenerator8x16[1570] = 8'he0;
assign _c_characterGenerator8x16[1571] = 8'h60;
assign _c_characterGenerator8x16[1572] = 8'h60;
assign _c_characterGenerator8x16[1573] = 8'h78;
assign _c_characterGenerator8x16[1574] = 8'h6c;
assign _c_characterGenerator8x16[1575] = 8'h66;
assign _c_characterGenerator8x16[1576] = 8'h66;
assign _c_characterGenerator8x16[1577] = 8'h66;
assign _c_characterGenerator8x16[1578] = 8'h66;
assign _c_characterGenerator8x16[1579] = 8'h7c;
assign _c_characterGenerator8x16[1580] = 8'h00;
assign _c_characterGenerator8x16[1581] = 8'h00;
assign _c_characterGenerator8x16[1582] = 8'h00;
assign _c_characterGenerator8x16[1583] = 8'h00;
assign _c_characterGenerator8x16[1584] = 8'h00;
assign _c_characterGenerator8x16[1585] = 8'h00;
assign _c_characterGenerator8x16[1586] = 8'h00;
assign _c_characterGenerator8x16[1587] = 8'h00;
assign _c_characterGenerator8x16[1588] = 8'h00;
assign _c_characterGenerator8x16[1589] = 8'h7c;
assign _c_characterGenerator8x16[1590] = 8'hc6;
assign _c_characterGenerator8x16[1591] = 8'hc0;
assign _c_characterGenerator8x16[1592] = 8'hc0;
assign _c_characterGenerator8x16[1593] = 8'hc0;
assign _c_characterGenerator8x16[1594] = 8'hc6;
assign _c_characterGenerator8x16[1595] = 8'h7c;
assign _c_characterGenerator8x16[1596] = 8'h00;
assign _c_characterGenerator8x16[1597] = 8'h00;
assign _c_characterGenerator8x16[1598] = 8'h00;
assign _c_characterGenerator8x16[1599] = 8'h00;
assign _c_characterGenerator8x16[1600] = 8'h00;
assign _c_characterGenerator8x16[1601] = 8'h00;
assign _c_characterGenerator8x16[1602] = 8'h1c;
assign _c_characterGenerator8x16[1603] = 8'h0c;
assign _c_characterGenerator8x16[1604] = 8'h0c;
assign _c_characterGenerator8x16[1605] = 8'h3c;
assign _c_characterGenerator8x16[1606] = 8'h6c;
assign _c_characterGenerator8x16[1607] = 8'hcc;
assign _c_characterGenerator8x16[1608] = 8'hcc;
assign _c_characterGenerator8x16[1609] = 8'hcc;
assign _c_characterGenerator8x16[1610] = 8'hcc;
assign _c_characterGenerator8x16[1611] = 8'h76;
assign _c_characterGenerator8x16[1612] = 8'h00;
assign _c_characterGenerator8x16[1613] = 8'h00;
assign _c_characterGenerator8x16[1614] = 8'h00;
assign _c_characterGenerator8x16[1615] = 8'h00;
assign _c_characterGenerator8x16[1616] = 8'h00;
assign _c_characterGenerator8x16[1617] = 8'h00;
assign _c_characterGenerator8x16[1618] = 8'h00;
assign _c_characterGenerator8x16[1619] = 8'h00;
assign _c_characterGenerator8x16[1620] = 8'h00;
assign _c_characterGenerator8x16[1621] = 8'h7c;
assign _c_characterGenerator8x16[1622] = 8'hc6;
assign _c_characterGenerator8x16[1623] = 8'hfe;
assign _c_characterGenerator8x16[1624] = 8'hc0;
assign _c_characterGenerator8x16[1625] = 8'hc0;
assign _c_characterGenerator8x16[1626] = 8'hc6;
assign _c_characterGenerator8x16[1627] = 8'h7c;
assign _c_characterGenerator8x16[1628] = 8'h00;
assign _c_characterGenerator8x16[1629] = 8'h00;
assign _c_characterGenerator8x16[1630] = 8'h00;
assign _c_characterGenerator8x16[1631] = 8'h00;
assign _c_characterGenerator8x16[1632] = 8'h00;
assign _c_characterGenerator8x16[1633] = 8'h00;
assign _c_characterGenerator8x16[1634] = 8'h38;
assign _c_characterGenerator8x16[1635] = 8'h6c;
assign _c_characterGenerator8x16[1636] = 8'h64;
assign _c_characterGenerator8x16[1637] = 8'h60;
assign _c_characterGenerator8x16[1638] = 8'hf0;
assign _c_characterGenerator8x16[1639] = 8'h60;
assign _c_characterGenerator8x16[1640] = 8'h60;
assign _c_characterGenerator8x16[1641] = 8'h60;
assign _c_characterGenerator8x16[1642] = 8'h60;
assign _c_characterGenerator8x16[1643] = 8'hf0;
assign _c_characterGenerator8x16[1644] = 8'h00;
assign _c_characterGenerator8x16[1645] = 8'h00;
assign _c_characterGenerator8x16[1646] = 8'h00;
assign _c_characterGenerator8x16[1647] = 8'h00;
assign _c_characterGenerator8x16[1648] = 8'h00;
assign _c_characterGenerator8x16[1649] = 8'h00;
assign _c_characterGenerator8x16[1650] = 8'h00;
assign _c_characterGenerator8x16[1651] = 8'h00;
assign _c_characterGenerator8x16[1652] = 8'h00;
assign _c_characterGenerator8x16[1653] = 8'h76;
assign _c_characterGenerator8x16[1654] = 8'hcc;
assign _c_characterGenerator8x16[1655] = 8'hcc;
assign _c_characterGenerator8x16[1656] = 8'hcc;
assign _c_characterGenerator8x16[1657] = 8'hcc;
assign _c_characterGenerator8x16[1658] = 8'hcc;
assign _c_characterGenerator8x16[1659] = 8'h7c;
assign _c_characterGenerator8x16[1660] = 8'h0c;
assign _c_characterGenerator8x16[1661] = 8'hcc;
assign _c_characterGenerator8x16[1662] = 8'h78;
assign _c_characterGenerator8x16[1663] = 8'h00;
assign _c_characterGenerator8x16[1664] = 8'h00;
assign _c_characterGenerator8x16[1665] = 8'h00;
assign _c_characterGenerator8x16[1666] = 8'he0;
assign _c_characterGenerator8x16[1667] = 8'h60;
assign _c_characterGenerator8x16[1668] = 8'h60;
assign _c_characterGenerator8x16[1669] = 8'h6c;
assign _c_characterGenerator8x16[1670] = 8'h76;
assign _c_characterGenerator8x16[1671] = 8'h66;
assign _c_characterGenerator8x16[1672] = 8'h66;
assign _c_characterGenerator8x16[1673] = 8'h66;
assign _c_characterGenerator8x16[1674] = 8'h66;
assign _c_characterGenerator8x16[1675] = 8'he6;
assign _c_characterGenerator8x16[1676] = 8'h00;
assign _c_characterGenerator8x16[1677] = 8'h00;
assign _c_characterGenerator8x16[1678] = 8'h00;
assign _c_characterGenerator8x16[1679] = 8'h00;
assign _c_characterGenerator8x16[1680] = 8'h00;
assign _c_characterGenerator8x16[1681] = 8'h00;
assign _c_characterGenerator8x16[1682] = 8'h18;
assign _c_characterGenerator8x16[1683] = 8'h18;
assign _c_characterGenerator8x16[1684] = 8'h00;
assign _c_characterGenerator8x16[1685] = 8'h38;
assign _c_characterGenerator8x16[1686] = 8'h18;
assign _c_characterGenerator8x16[1687] = 8'h18;
assign _c_characterGenerator8x16[1688] = 8'h18;
assign _c_characterGenerator8x16[1689] = 8'h18;
assign _c_characterGenerator8x16[1690] = 8'h18;
assign _c_characterGenerator8x16[1691] = 8'h3c;
assign _c_characterGenerator8x16[1692] = 8'h00;
assign _c_characterGenerator8x16[1693] = 8'h00;
assign _c_characterGenerator8x16[1694] = 8'h00;
assign _c_characterGenerator8x16[1695] = 8'h00;
assign _c_characterGenerator8x16[1696] = 8'h00;
assign _c_characterGenerator8x16[1697] = 8'h00;
assign _c_characterGenerator8x16[1698] = 8'h06;
assign _c_characterGenerator8x16[1699] = 8'h06;
assign _c_characterGenerator8x16[1700] = 8'h00;
assign _c_characterGenerator8x16[1701] = 8'h0e;
assign _c_characterGenerator8x16[1702] = 8'h06;
assign _c_characterGenerator8x16[1703] = 8'h06;
assign _c_characterGenerator8x16[1704] = 8'h06;
assign _c_characterGenerator8x16[1705] = 8'h06;
assign _c_characterGenerator8x16[1706] = 8'h06;
assign _c_characterGenerator8x16[1707] = 8'h06;
assign _c_characterGenerator8x16[1708] = 8'h66;
assign _c_characterGenerator8x16[1709] = 8'h66;
assign _c_characterGenerator8x16[1710] = 8'h3c;
assign _c_characterGenerator8x16[1711] = 8'h00;
assign _c_characterGenerator8x16[1712] = 8'h00;
assign _c_characterGenerator8x16[1713] = 8'h00;
assign _c_characterGenerator8x16[1714] = 8'he0;
assign _c_characterGenerator8x16[1715] = 8'h60;
assign _c_characterGenerator8x16[1716] = 8'h60;
assign _c_characterGenerator8x16[1717] = 8'h66;
assign _c_characterGenerator8x16[1718] = 8'h6c;
assign _c_characterGenerator8x16[1719] = 8'h78;
assign _c_characterGenerator8x16[1720] = 8'h78;
assign _c_characterGenerator8x16[1721] = 8'h6c;
assign _c_characterGenerator8x16[1722] = 8'h66;
assign _c_characterGenerator8x16[1723] = 8'he6;
assign _c_characterGenerator8x16[1724] = 8'h00;
assign _c_characterGenerator8x16[1725] = 8'h00;
assign _c_characterGenerator8x16[1726] = 8'h00;
assign _c_characterGenerator8x16[1727] = 8'h00;
assign _c_characterGenerator8x16[1728] = 8'h00;
assign _c_characterGenerator8x16[1729] = 8'h00;
assign _c_characterGenerator8x16[1730] = 8'h38;
assign _c_characterGenerator8x16[1731] = 8'h18;
assign _c_characterGenerator8x16[1732] = 8'h18;
assign _c_characterGenerator8x16[1733] = 8'h18;
assign _c_characterGenerator8x16[1734] = 8'h18;
assign _c_characterGenerator8x16[1735] = 8'h18;
assign _c_characterGenerator8x16[1736] = 8'h18;
assign _c_characterGenerator8x16[1737] = 8'h18;
assign _c_characterGenerator8x16[1738] = 8'h18;
assign _c_characterGenerator8x16[1739] = 8'h3c;
assign _c_characterGenerator8x16[1740] = 8'h00;
assign _c_characterGenerator8x16[1741] = 8'h00;
assign _c_characterGenerator8x16[1742] = 8'h00;
assign _c_characterGenerator8x16[1743] = 8'h00;
assign _c_characterGenerator8x16[1744] = 8'h00;
assign _c_characterGenerator8x16[1745] = 8'h00;
assign _c_characterGenerator8x16[1746] = 8'h00;
assign _c_characterGenerator8x16[1747] = 8'h00;
assign _c_characterGenerator8x16[1748] = 8'h00;
assign _c_characterGenerator8x16[1749] = 8'hec;
assign _c_characterGenerator8x16[1750] = 8'hfe;
assign _c_characterGenerator8x16[1751] = 8'hd6;
assign _c_characterGenerator8x16[1752] = 8'hd6;
assign _c_characterGenerator8x16[1753] = 8'hd6;
assign _c_characterGenerator8x16[1754] = 8'hd6;
assign _c_characterGenerator8x16[1755] = 8'hc6;
assign _c_characterGenerator8x16[1756] = 8'h00;
assign _c_characterGenerator8x16[1757] = 8'h00;
assign _c_characterGenerator8x16[1758] = 8'h00;
assign _c_characterGenerator8x16[1759] = 8'h00;
assign _c_characterGenerator8x16[1760] = 8'h00;
assign _c_characterGenerator8x16[1761] = 8'h00;
assign _c_characterGenerator8x16[1762] = 8'h00;
assign _c_characterGenerator8x16[1763] = 8'h00;
assign _c_characterGenerator8x16[1764] = 8'h00;
assign _c_characterGenerator8x16[1765] = 8'hdc;
assign _c_characterGenerator8x16[1766] = 8'h66;
assign _c_characterGenerator8x16[1767] = 8'h66;
assign _c_characterGenerator8x16[1768] = 8'h66;
assign _c_characterGenerator8x16[1769] = 8'h66;
assign _c_characterGenerator8x16[1770] = 8'h66;
assign _c_characterGenerator8x16[1771] = 8'h66;
assign _c_characterGenerator8x16[1772] = 8'h00;
assign _c_characterGenerator8x16[1773] = 8'h00;
assign _c_characterGenerator8x16[1774] = 8'h00;
assign _c_characterGenerator8x16[1775] = 8'h00;
assign _c_characterGenerator8x16[1776] = 8'h00;
assign _c_characterGenerator8x16[1777] = 8'h00;
assign _c_characterGenerator8x16[1778] = 8'h00;
assign _c_characterGenerator8x16[1779] = 8'h00;
assign _c_characterGenerator8x16[1780] = 8'h00;
assign _c_characterGenerator8x16[1781] = 8'h7c;
assign _c_characterGenerator8x16[1782] = 8'hc6;
assign _c_characterGenerator8x16[1783] = 8'hc6;
assign _c_characterGenerator8x16[1784] = 8'hc6;
assign _c_characterGenerator8x16[1785] = 8'hc6;
assign _c_characterGenerator8x16[1786] = 8'hc6;
assign _c_characterGenerator8x16[1787] = 8'h7c;
assign _c_characterGenerator8x16[1788] = 8'h00;
assign _c_characterGenerator8x16[1789] = 8'h00;
assign _c_characterGenerator8x16[1790] = 8'h00;
assign _c_characterGenerator8x16[1791] = 8'h00;
assign _c_characterGenerator8x16[1792] = 8'h00;
assign _c_characterGenerator8x16[1793] = 8'h00;
assign _c_characterGenerator8x16[1794] = 8'h00;
assign _c_characterGenerator8x16[1795] = 8'h00;
assign _c_characterGenerator8x16[1796] = 8'h00;
assign _c_characterGenerator8x16[1797] = 8'hdc;
assign _c_characterGenerator8x16[1798] = 8'h66;
assign _c_characterGenerator8x16[1799] = 8'h66;
assign _c_characterGenerator8x16[1800] = 8'h66;
assign _c_characterGenerator8x16[1801] = 8'h66;
assign _c_characterGenerator8x16[1802] = 8'h66;
assign _c_characterGenerator8x16[1803] = 8'h7c;
assign _c_characterGenerator8x16[1804] = 8'h60;
assign _c_characterGenerator8x16[1805] = 8'h60;
assign _c_characterGenerator8x16[1806] = 8'hf0;
assign _c_characterGenerator8x16[1807] = 8'h00;
assign _c_characterGenerator8x16[1808] = 8'h00;
assign _c_characterGenerator8x16[1809] = 8'h00;
assign _c_characterGenerator8x16[1810] = 8'h00;
assign _c_characterGenerator8x16[1811] = 8'h00;
assign _c_characterGenerator8x16[1812] = 8'h00;
assign _c_characterGenerator8x16[1813] = 8'h76;
assign _c_characterGenerator8x16[1814] = 8'hcc;
assign _c_characterGenerator8x16[1815] = 8'hcc;
assign _c_characterGenerator8x16[1816] = 8'hcc;
assign _c_characterGenerator8x16[1817] = 8'hcc;
assign _c_characterGenerator8x16[1818] = 8'hcc;
assign _c_characterGenerator8x16[1819] = 8'h7c;
assign _c_characterGenerator8x16[1820] = 8'h0c;
assign _c_characterGenerator8x16[1821] = 8'h0c;
assign _c_characterGenerator8x16[1822] = 8'h1e;
assign _c_characterGenerator8x16[1823] = 8'h00;
assign _c_characterGenerator8x16[1824] = 8'h00;
assign _c_characterGenerator8x16[1825] = 8'h00;
assign _c_characterGenerator8x16[1826] = 8'h00;
assign _c_characterGenerator8x16[1827] = 8'h00;
assign _c_characterGenerator8x16[1828] = 8'h00;
assign _c_characterGenerator8x16[1829] = 8'hdc;
assign _c_characterGenerator8x16[1830] = 8'h76;
assign _c_characterGenerator8x16[1831] = 8'h66;
assign _c_characterGenerator8x16[1832] = 8'h60;
assign _c_characterGenerator8x16[1833] = 8'h60;
assign _c_characterGenerator8x16[1834] = 8'h60;
assign _c_characterGenerator8x16[1835] = 8'hf0;
assign _c_characterGenerator8x16[1836] = 8'h00;
assign _c_characterGenerator8x16[1837] = 8'h00;
assign _c_characterGenerator8x16[1838] = 8'h00;
assign _c_characterGenerator8x16[1839] = 8'h00;
assign _c_characterGenerator8x16[1840] = 8'h00;
assign _c_characterGenerator8x16[1841] = 8'h00;
assign _c_characterGenerator8x16[1842] = 8'h00;
assign _c_characterGenerator8x16[1843] = 8'h00;
assign _c_characterGenerator8x16[1844] = 8'h00;
assign _c_characterGenerator8x16[1845] = 8'h7c;
assign _c_characterGenerator8x16[1846] = 8'hc6;
assign _c_characterGenerator8x16[1847] = 8'h60;
assign _c_characterGenerator8x16[1848] = 8'h38;
assign _c_characterGenerator8x16[1849] = 8'h0c;
assign _c_characterGenerator8x16[1850] = 8'hc6;
assign _c_characterGenerator8x16[1851] = 8'h7c;
assign _c_characterGenerator8x16[1852] = 8'h00;
assign _c_characterGenerator8x16[1853] = 8'h00;
assign _c_characterGenerator8x16[1854] = 8'h00;
assign _c_characterGenerator8x16[1855] = 8'h00;
assign _c_characterGenerator8x16[1856] = 8'h00;
assign _c_characterGenerator8x16[1857] = 8'h00;
assign _c_characterGenerator8x16[1858] = 8'h10;
assign _c_characterGenerator8x16[1859] = 8'h30;
assign _c_characterGenerator8x16[1860] = 8'h30;
assign _c_characterGenerator8x16[1861] = 8'hfc;
assign _c_characterGenerator8x16[1862] = 8'h30;
assign _c_characterGenerator8x16[1863] = 8'h30;
assign _c_characterGenerator8x16[1864] = 8'h30;
assign _c_characterGenerator8x16[1865] = 8'h30;
assign _c_characterGenerator8x16[1866] = 8'h36;
assign _c_characterGenerator8x16[1867] = 8'h1c;
assign _c_characterGenerator8x16[1868] = 8'h00;
assign _c_characterGenerator8x16[1869] = 8'h00;
assign _c_characterGenerator8x16[1870] = 8'h00;
assign _c_characterGenerator8x16[1871] = 8'h00;
assign _c_characterGenerator8x16[1872] = 8'h00;
assign _c_characterGenerator8x16[1873] = 8'h00;
assign _c_characterGenerator8x16[1874] = 8'h00;
assign _c_characterGenerator8x16[1875] = 8'h00;
assign _c_characterGenerator8x16[1876] = 8'h00;
assign _c_characterGenerator8x16[1877] = 8'hcc;
assign _c_characterGenerator8x16[1878] = 8'hcc;
assign _c_characterGenerator8x16[1879] = 8'hcc;
assign _c_characterGenerator8x16[1880] = 8'hcc;
assign _c_characterGenerator8x16[1881] = 8'hcc;
assign _c_characterGenerator8x16[1882] = 8'hcc;
assign _c_characterGenerator8x16[1883] = 8'h76;
assign _c_characterGenerator8x16[1884] = 8'h00;
assign _c_characterGenerator8x16[1885] = 8'h00;
assign _c_characterGenerator8x16[1886] = 8'h00;
assign _c_characterGenerator8x16[1887] = 8'h00;
assign _c_characterGenerator8x16[1888] = 8'h00;
assign _c_characterGenerator8x16[1889] = 8'h00;
assign _c_characterGenerator8x16[1890] = 8'h00;
assign _c_characterGenerator8x16[1891] = 8'h00;
assign _c_characterGenerator8x16[1892] = 8'h00;
assign _c_characterGenerator8x16[1893] = 8'h66;
assign _c_characterGenerator8x16[1894] = 8'h66;
assign _c_characterGenerator8x16[1895] = 8'h66;
assign _c_characterGenerator8x16[1896] = 8'h66;
assign _c_characterGenerator8x16[1897] = 8'h66;
assign _c_characterGenerator8x16[1898] = 8'h3c;
assign _c_characterGenerator8x16[1899] = 8'h18;
assign _c_characterGenerator8x16[1900] = 8'h00;
assign _c_characterGenerator8x16[1901] = 8'h00;
assign _c_characterGenerator8x16[1902] = 8'h00;
assign _c_characterGenerator8x16[1903] = 8'h00;
assign _c_characterGenerator8x16[1904] = 8'h00;
assign _c_characterGenerator8x16[1905] = 8'h00;
assign _c_characterGenerator8x16[1906] = 8'h00;
assign _c_characterGenerator8x16[1907] = 8'h00;
assign _c_characterGenerator8x16[1908] = 8'h00;
assign _c_characterGenerator8x16[1909] = 8'hc6;
assign _c_characterGenerator8x16[1910] = 8'hc6;
assign _c_characterGenerator8x16[1911] = 8'hd6;
assign _c_characterGenerator8x16[1912] = 8'hd6;
assign _c_characterGenerator8x16[1913] = 8'hd6;
assign _c_characterGenerator8x16[1914] = 8'hfe;
assign _c_characterGenerator8x16[1915] = 8'h6c;
assign _c_characterGenerator8x16[1916] = 8'h00;
assign _c_characterGenerator8x16[1917] = 8'h00;
assign _c_characterGenerator8x16[1918] = 8'h00;
assign _c_characterGenerator8x16[1919] = 8'h00;
assign _c_characterGenerator8x16[1920] = 8'h00;
assign _c_characterGenerator8x16[1921] = 8'h00;
assign _c_characterGenerator8x16[1922] = 8'h00;
assign _c_characterGenerator8x16[1923] = 8'h00;
assign _c_characterGenerator8x16[1924] = 8'h00;
assign _c_characterGenerator8x16[1925] = 8'hc6;
assign _c_characterGenerator8x16[1926] = 8'h6c;
assign _c_characterGenerator8x16[1927] = 8'h38;
assign _c_characterGenerator8x16[1928] = 8'h38;
assign _c_characterGenerator8x16[1929] = 8'h38;
assign _c_characterGenerator8x16[1930] = 8'h6c;
assign _c_characterGenerator8x16[1931] = 8'hc6;
assign _c_characterGenerator8x16[1932] = 8'h00;
assign _c_characterGenerator8x16[1933] = 8'h00;
assign _c_characterGenerator8x16[1934] = 8'h00;
assign _c_characterGenerator8x16[1935] = 8'h00;
assign _c_characterGenerator8x16[1936] = 8'h00;
assign _c_characterGenerator8x16[1937] = 8'h00;
assign _c_characterGenerator8x16[1938] = 8'h00;
assign _c_characterGenerator8x16[1939] = 8'h00;
assign _c_characterGenerator8x16[1940] = 8'h00;
assign _c_characterGenerator8x16[1941] = 8'hc6;
assign _c_characterGenerator8x16[1942] = 8'hc6;
assign _c_characterGenerator8x16[1943] = 8'hc6;
assign _c_characterGenerator8x16[1944] = 8'hc6;
assign _c_characterGenerator8x16[1945] = 8'hc6;
assign _c_characterGenerator8x16[1946] = 8'hc6;
assign _c_characterGenerator8x16[1947] = 8'h7e;
assign _c_characterGenerator8x16[1948] = 8'h06;
assign _c_characterGenerator8x16[1949] = 8'h0c;
assign _c_characterGenerator8x16[1950] = 8'hf8;
assign _c_characterGenerator8x16[1951] = 8'h00;
assign _c_characterGenerator8x16[1952] = 8'h00;
assign _c_characterGenerator8x16[1953] = 8'h00;
assign _c_characterGenerator8x16[1954] = 8'h00;
assign _c_characterGenerator8x16[1955] = 8'h00;
assign _c_characterGenerator8x16[1956] = 8'h00;
assign _c_characterGenerator8x16[1957] = 8'hfe;
assign _c_characterGenerator8x16[1958] = 8'hcc;
assign _c_characterGenerator8x16[1959] = 8'h18;
assign _c_characterGenerator8x16[1960] = 8'h30;
assign _c_characterGenerator8x16[1961] = 8'h60;
assign _c_characterGenerator8x16[1962] = 8'hc6;
assign _c_characterGenerator8x16[1963] = 8'hfe;
assign _c_characterGenerator8x16[1964] = 8'h00;
assign _c_characterGenerator8x16[1965] = 8'h00;
assign _c_characterGenerator8x16[1966] = 8'h00;
assign _c_characterGenerator8x16[1967] = 8'h00;
assign _c_characterGenerator8x16[1968] = 8'h00;
assign _c_characterGenerator8x16[1969] = 8'h00;
assign _c_characterGenerator8x16[1970] = 8'h0e;
assign _c_characterGenerator8x16[1971] = 8'h18;
assign _c_characterGenerator8x16[1972] = 8'h18;
assign _c_characterGenerator8x16[1973] = 8'h18;
assign _c_characterGenerator8x16[1974] = 8'h70;
assign _c_characterGenerator8x16[1975] = 8'h18;
assign _c_characterGenerator8x16[1976] = 8'h18;
assign _c_characterGenerator8x16[1977] = 8'h18;
assign _c_characterGenerator8x16[1978] = 8'h18;
assign _c_characterGenerator8x16[1979] = 8'h0e;
assign _c_characterGenerator8x16[1980] = 8'h00;
assign _c_characterGenerator8x16[1981] = 8'h00;
assign _c_characterGenerator8x16[1982] = 8'h00;
assign _c_characterGenerator8x16[1983] = 8'h00;
assign _c_characterGenerator8x16[1984] = 8'h00;
assign _c_characterGenerator8x16[1985] = 8'h00;
assign _c_characterGenerator8x16[1986] = 8'h18;
assign _c_characterGenerator8x16[1987] = 8'h18;
assign _c_characterGenerator8x16[1988] = 8'h18;
assign _c_characterGenerator8x16[1989] = 8'h18;
assign _c_characterGenerator8x16[1990] = 8'h00;
assign _c_characterGenerator8x16[1991] = 8'h18;
assign _c_characterGenerator8x16[1992] = 8'h18;
assign _c_characterGenerator8x16[1993] = 8'h18;
assign _c_characterGenerator8x16[1994] = 8'h18;
assign _c_characterGenerator8x16[1995] = 8'h18;
assign _c_characterGenerator8x16[1996] = 8'h00;
assign _c_characterGenerator8x16[1997] = 8'h00;
assign _c_characterGenerator8x16[1998] = 8'h00;
assign _c_characterGenerator8x16[1999] = 8'h00;
assign _c_characterGenerator8x16[2000] = 8'h00;
assign _c_characterGenerator8x16[2001] = 8'h00;
assign _c_characterGenerator8x16[2002] = 8'h70;
assign _c_characterGenerator8x16[2003] = 8'h18;
assign _c_characterGenerator8x16[2004] = 8'h18;
assign _c_characterGenerator8x16[2005] = 8'h18;
assign _c_characterGenerator8x16[2006] = 8'h0e;
assign _c_characterGenerator8x16[2007] = 8'h18;
assign _c_characterGenerator8x16[2008] = 8'h18;
assign _c_characterGenerator8x16[2009] = 8'h18;
assign _c_characterGenerator8x16[2010] = 8'h18;
assign _c_characterGenerator8x16[2011] = 8'h70;
assign _c_characterGenerator8x16[2012] = 8'h00;
assign _c_characterGenerator8x16[2013] = 8'h00;
assign _c_characterGenerator8x16[2014] = 8'h00;
assign _c_characterGenerator8x16[2015] = 8'h00;
assign _c_characterGenerator8x16[2016] = 8'h00;
assign _c_characterGenerator8x16[2017] = 8'h00;
assign _c_characterGenerator8x16[2018] = 8'h76;
assign _c_characterGenerator8x16[2019] = 8'hdc;
assign _c_characterGenerator8x16[2020] = 8'h00;
assign _c_characterGenerator8x16[2021] = 8'h00;
assign _c_characterGenerator8x16[2022] = 8'h00;
assign _c_characterGenerator8x16[2023] = 8'h00;
assign _c_characterGenerator8x16[2024] = 8'h00;
assign _c_characterGenerator8x16[2025] = 8'h00;
assign _c_characterGenerator8x16[2026] = 8'h00;
assign _c_characterGenerator8x16[2027] = 8'h00;
assign _c_characterGenerator8x16[2028] = 8'h00;
assign _c_characterGenerator8x16[2029] = 8'h00;
assign _c_characterGenerator8x16[2030] = 8'h00;
assign _c_characterGenerator8x16[2031] = 8'h00;
assign _c_characterGenerator8x16[2032] = 8'h00;
assign _c_characterGenerator8x16[2033] = 8'h00;
assign _c_characterGenerator8x16[2034] = 8'h00;
assign _c_characterGenerator8x16[2035] = 8'h00;
assign _c_characterGenerator8x16[2036] = 8'h10;
assign _c_characterGenerator8x16[2037] = 8'h38;
assign _c_characterGenerator8x16[2038] = 8'h6c;
assign _c_characterGenerator8x16[2039] = 8'hc6;
assign _c_characterGenerator8x16[2040] = 8'hc6;
assign _c_characterGenerator8x16[2041] = 8'hc6;
assign _c_characterGenerator8x16[2042] = 8'hfe;
assign _c_characterGenerator8x16[2043] = 8'h00;
assign _c_characterGenerator8x16[2044] = 8'h00;
assign _c_characterGenerator8x16[2045] = 8'h00;
assign _c_characterGenerator8x16[2046] = 8'h00;
assign _c_characterGenerator8x16[2047] = 8'h00;
assign _c_characterGenerator8x16[2048] = 8'h00;
assign _c_characterGenerator8x16[2049] = 8'h00;
assign _c_characterGenerator8x16[2050] = 8'h3c;
assign _c_characterGenerator8x16[2051] = 8'h66;
assign _c_characterGenerator8x16[2052] = 8'hc2;
assign _c_characterGenerator8x16[2053] = 8'hc0;
assign _c_characterGenerator8x16[2054] = 8'hc0;
assign _c_characterGenerator8x16[2055] = 8'hc0;
assign _c_characterGenerator8x16[2056] = 8'hc2;
assign _c_characterGenerator8x16[2057] = 8'h66;
assign _c_characterGenerator8x16[2058] = 8'h3c;
assign _c_characterGenerator8x16[2059] = 8'h0c;
assign _c_characterGenerator8x16[2060] = 8'h06;
assign _c_characterGenerator8x16[2061] = 8'h7c;
assign _c_characterGenerator8x16[2062] = 8'h00;
assign _c_characterGenerator8x16[2063] = 8'h00;
assign _c_characterGenerator8x16[2064] = 8'h00;
assign _c_characterGenerator8x16[2065] = 8'h00;
assign _c_characterGenerator8x16[2066] = 8'hcc;
assign _c_characterGenerator8x16[2067] = 8'h00;
assign _c_characterGenerator8x16[2068] = 8'h00;
assign _c_characterGenerator8x16[2069] = 8'hcc;
assign _c_characterGenerator8x16[2070] = 8'hcc;
assign _c_characterGenerator8x16[2071] = 8'hcc;
assign _c_characterGenerator8x16[2072] = 8'hcc;
assign _c_characterGenerator8x16[2073] = 8'hcc;
assign _c_characterGenerator8x16[2074] = 8'hcc;
assign _c_characterGenerator8x16[2075] = 8'h76;
assign _c_characterGenerator8x16[2076] = 8'h00;
assign _c_characterGenerator8x16[2077] = 8'h00;
assign _c_characterGenerator8x16[2078] = 8'h00;
assign _c_characterGenerator8x16[2079] = 8'h00;
assign _c_characterGenerator8x16[2080] = 8'h00;
assign _c_characterGenerator8x16[2081] = 8'h0c;
assign _c_characterGenerator8x16[2082] = 8'h18;
assign _c_characterGenerator8x16[2083] = 8'h30;
assign _c_characterGenerator8x16[2084] = 8'h00;
assign _c_characterGenerator8x16[2085] = 8'h7c;
assign _c_characterGenerator8x16[2086] = 8'hc6;
assign _c_characterGenerator8x16[2087] = 8'hfe;
assign _c_characterGenerator8x16[2088] = 8'hc0;
assign _c_characterGenerator8x16[2089] = 8'hc0;
assign _c_characterGenerator8x16[2090] = 8'hc6;
assign _c_characterGenerator8x16[2091] = 8'h7c;
assign _c_characterGenerator8x16[2092] = 8'h00;
assign _c_characterGenerator8x16[2093] = 8'h00;
assign _c_characterGenerator8x16[2094] = 8'h00;
assign _c_characterGenerator8x16[2095] = 8'h00;
assign _c_characterGenerator8x16[2096] = 8'h00;
assign _c_characterGenerator8x16[2097] = 8'h10;
assign _c_characterGenerator8x16[2098] = 8'h38;
assign _c_characterGenerator8x16[2099] = 8'h6c;
assign _c_characterGenerator8x16[2100] = 8'h00;
assign _c_characterGenerator8x16[2101] = 8'h78;
assign _c_characterGenerator8x16[2102] = 8'h0c;
assign _c_characterGenerator8x16[2103] = 8'h7c;
assign _c_characterGenerator8x16[2104] = 8'hcc;
assign _c_characterGenerator8x16[2105] = 8'hcc;
assign _c_characterGenerator8x16[2106] = 8'hcc;
assign _c_characterGenerator8x16[2107] = 8'h76;
assign _c_characterGenerator8x16[2108] = 8'h00;
assign _c_characterGenerator8x16[2109] = 8'h00;
assign _c_characterGenerator8x16[2110] = 8'h00;
assign _c_characterGenerator8x16[2111] = 8'h00;
assign _c_characterGenerator8x16[2112] = 8'h00;
assign _c_characterGenerator8x16[2113] = 8'h00;
assign _c_characterGenerator8x16[2114] = 8'hcc;
assign _c_characterGenerator8x16[2115] = 8'h00;
assign _c_characterGenerator8x16[2116] = 8'h00;
assign _c_characterGenerator8x16[2117] = 8'h78;
assign _c_characterGenerator8x16[2118] = 8'h0c;
assign _c_characterGenerator8x16[2119] = 8'h7c;
assign _c_characterGenerator8x16[2120] = 8'hcc;
assign _c_characterGenerator8x16[2121] = 8'hcc;
assign _c_characterGenerator8x16[2122] = 8'hcc;
assign _c_characterGenerator8x16[2123] = 8'h76;
assign _c_characterGenerator8x16[2124] = 8'h00;
assign _c_characterGenerator8x16[2125] = 8'h00;
assign _c_characterGenerator8x16[2126] = 8'h00;
assign _c_characterGenerator8x16[2127] = 8'h00;
assign _c_characterGenerator8x16[2128] = 8'h00;
assign _c_characterGenerator8x16[2129] = 8'h60;
assign _c_characterGenerator8x16[2130] = 8'h30;
assign _c_characterGenerator8x16[2131] = 8'h18;
assign _c_characterGenerator8x16[2132] = 8'h00;
assign _c_characterGenerator8x16[2133] = 8'h78;
assign _c_characterGenerator8x16[2134] = 8'h0c;
assign _c_characterGenerator8x16[2135] = 8'h7c;
assign _c_characterGenerator8x16[2136] = 8'hcc;
assign _c_characterGenerator8x16[2137] = 8'hcc;
assign _c_characterGenerator8x16[2138] = 8'hcc;
assign _c_characterGenerator8x16[2139] = 8'h76;
assign _c_characterGenerator8x16[2140] = 8'h00;
assign _c_characterGenerator8x16[2141] = 8'h00;
assign _c_characterGenerator8x16[2142] = 8'h00;
assign _c_characterGenerator8x16[2143] = 8'h00;
assign _c_characterGenerator8x16[2144] = 8'h00;
assign _c_characterGenerator8x16[2145] = 8'h38;
assign _c_characterGenerator8x16[2146] = 8'h6c;
assign _c_characterGenerator8x16[2147] = 8'h38;
assign _c_characterGenerator8x16[2148] = 8'h00;
assign _c_characterGenerator8x16[2149] = 8'h78;
assign _c_characterGenerator8x16[2150] = 8'h0c;
assign _c_characterGenerator8x16[2151] = 8'h7c;
assign _c_characterGenerator8x16[2152] = 8'hcc;
assign _c_characterGenerator8x16[2153] = 8'hcc;
assign _c_characterGenerator8x16[2154] = 8'hcc;
assign _c_characterGenerator8x16[2155] = 8'h76;
assign _c_characterGenerator8x16[2156] = 8'h00;
assign _c_characterGenerator8x16[2157] = 8'h00;
assign _c_characterGenerator8x16[2158] = 8'h00;
assign _c_characterGenerator8x16[2159] = 8'h00;
assign _c_characterGenerator8x16[2160] = 8'h00;
assign _c_characterGenerator8x16[2161] = 8'h00;
assign _c_characterGenerator8x16[2162] = 8'h00;
assign _c_characterGenerator8x16[2163] = 8'h00;
assign _c_characterGenerator8x16[2164] = 8'h3c;
assign _c_characterGenerator8x16[2165] = 8'h66;
assign _c_characterGenerator8x16[2166] = 8'h60;
assign _c_characterGenerator8x16[2167] = 8'h60;
assign _c_characterGenerator8x16[2168] = 8'h66;
assign _c_characterGenerator8x16[2169] = 8'h3c;
assign _c_characterGenerator8x16[2170] = 8'h0c;
assign _c_characterGenerator8x16[2171] = 8'h06;
assign _c_characterGenerator8x16[2172] = 8'h3c;
assign _c_characterGenerator8x16[2173] = 8'h00;
assign _c_characterGenerator8x16[2174] = 8'h00;
assign _c_characterGenerator8x16[2175] = 8'h00;
assign _c_characterGenerator8x16[2176] = 8'h00;
assign _c_characterGenerator8x16[2177] = 8'h10;
assign _c_characterGenerator8x16[2178] = 8'h38;
assign _c_characterGenerator8x16[2179] = 8'h6c;
assign _c_characterGenerator8x16[2180] = 8'h00;
assign _c_characterGenerator8x16[2181] = 8'h7c;
assign _c_characterGenerator8x16[2182] = 8'hc6;
assign _c_characterGenerator8x16[2183] = 8'hfe;
assign _c_characterGenerator8x16[2184] = 8'hc0;
assign _c_characterGenerator8x16[2185] = 8'hc0;
assign _c_characterGenerator8x16[2186] = 8'hc6;
assign _c_characterGenerator8x16[2187] = 8'h7c;
assign _c_characterGenerator8x16[2188] = 8'h00;
assign _c_characterGenerator8x16[2189] = 8'h00;
assign _c_characterGenerator8x16[2190] = 8'h00;
assign _c_characterGenerator8x16[2191] = 8'h00;
assign _c_characterGenerator8x16[2192] = 8'h00;
assign _c_characterGenerator8x16[2193] = 8'h00;
assign _c_characterGenerator8x16[2194] = 8'hc6;
assign _c_characterGenerator8x16[2195] = 8'h00;
assign _c_characterGenerator8x16[2196] = 8'h00;
assign _c_characterGenerator8x16[2197] = 8'h7c;
assign _c_characterGenerator8x16[2198] = 8'hc6;
assign _c_characterGenerator8x16[2199] = 8'hfe;
assign _c_characterGenerator8x16[2200] = 8'hc0;
assign _c_characterGenerator8x16[2201] = 8'hc0;
assign _c_characterGenerator8x16[2202] = 8'hc6;
assign _c_characterGenerator8x16[2203] = 8'h7c;
assign _c_characterGenerator8x16[2204] = 8'h00;
assign _c_characterGenerator8x16[2205] = 8'h00;
assign _c_characterGenerator8x16[2206] = 8'h00;
assign _c_characterGenerator8x16[2207] = 8'h00;
assign _c_characterGenerator8x16[2208] = 8'h00;
assign _c_characterGenerator8x16[2209] = 8'h60;
assign _c_characterGenerator8x16[2210] = 8'h30;
assign _c_characterGenerator8x16[2211] = 8'h18;
assign _c_characterGenerator8x16[2212] = 8'h00;
assign _c_characterGenerator8x16[2213] = 8'h7c;
assign _c_characterGenerator8x16[2214] = 8'hc6;
assign _c_characterGenerator8x16[2215] = 8'hfe;
assign _c_characterGenerator8x16[2216] = 8'hc0;
assign _c_characterGenerator8x16[2217] = 8'hc0;
assign _c_characterGenerator8x16[2218] = 8'hc6;
assign _c_characterGenerator8x16[2219] = 8'h7c;
assign _c_characterGenerator8x16[2220] = 8'h00;
assign _c_characterGenerator8x16[2221] = 8'h00;
assign _c_characterGenerator8x16[2222] = 8'h00;
assign _c_characterGenerator8x16[2223] = 8'h00;
assign _c_characterGenerator8x16[2224] = 8'h00;
assign _c_characterGenerator8x16[2225] = 8'h00;
assign _c_characterGenerator8x16[2226] = 8'h66;
assign _c_characterGenerator8x16[2227] = 8'h00;
assign _c_characterGenerator8x16[2228] = 8'h00;
assign _c_characterGenerator8x16[2229] = 8'h38;
assign _c_characterGenerator8x16[2230] = 8'h18;
assign _c_characterGenerator8x16[2231] = 8'h18;
assign _c_characterGenerator8x16[2232] = 8'h18;
assign _c_characterGenerator8x16[2233] = 8'h18;
assign _c_characterGenerator8x16[2234] = 8'h18;
assign _c_characterGenerator8x16[2235] = 8'h3c;
assign _c_characterGenerator8x16[2236] = 8'h00;
assign _c_characterGenerator8x16[2237] = 8'h00;
assign _c_characterGenerator8x16[2238] = 8'h00;
assign _c_characterGenerator8x16[2239] = 8'h00;
assign _c_characterGenerator8x16[2240] = 8'h00;
assign _c_characterGenerator8x16[2241] = 8'h18;
assign _c_characterGenerator8x16[2242] = 8'h3c;
assign _c_characterGenerator8x16[2243] = 8'h66;
assign _c_characterGenerator8x16[2244] = 8'h00;
assign _c_characterGenerator8x16[2245] = 8'h38;
assign _c_characterGenerator8x16[2246] = 8'h18;
assign _c_characterGenerator8x16[2247] = 8'h18;
assign _c_characterGenerator8x16[2248] = 8'h18;
assign _c_characterGenerator8x16[2249] = 8'h18;
assign _c_characterGenerator8x16[2250] = 8'h18;
assign _c_characterGenerator8x16[2251] = 8'h3c;
assign _c_characterGenerator8x16[2252] = 8'h00;
assign _c_characterGenerator8x16[2253] = 8'h00;
assign _c_characterGenerator8x16[2254] = 8'h00;
assign _c_characterGenerator8x16[2255] = 8'h00;
assign _c_characterGenerator8x16[2256] = 8'h00;
assign _c_characterGenerator8x16[2257] = 8'h60;
assign _c_characterGenerator8x16[2258] = 8'h30;
assign _c_characterGenerator8x16[2259] = 8'h18;
assign _c_characterGenerator8x16[2260] = 8'h00;
assign _c_characterGenerator8x16[2261] = 8'h38;
assign _c_characterGenerator8x16[2262] = 8'h18;
assign _c_characterGenerator8x16[2263] = 8'h18;
assign _c_characterGenerator8x16[2264] = 8'h18;
assign _c_characterGenerator8x16[2265] = 8'h18;
assign _c_characterGenerator8x16[2266] = 8'h18;
assign _c_characterGenerator8x16[2267] = 8'h3c;
assign _c_characterGenerator8x16[2268] = 8'h00;
assign _c_characterGenerator8x16[2269] = 8'h00;
assign _c_characterGenerator8x16[2270] = 8'h00;
assign _c_characterGenerator8x16[2271] = 8'h00;
assign _c_characterGenerator8x16[2272] = 8'h00;
assign _c_characterGenerator8x16[2273] = 8'hc6;
assign _c_characterGenerator8x16[2274] = 8'h00;
assign _c_characterGenerator8x16[2275] = 8'h10;
assign _c_characterGenerator8x16[2276] = 8'h38;
assign _c_characterGenerator8x16[2277] = 8'h6c;
assign _c_characterGenerator8x16[2278] = 8'hc6;
assign _c_characterGenerator8x16[2279] = 8'hc6;
assign _c_characterGenerator8x16[2280] = 8'hfe;
assign _c_characterGenerator8x16[2281] = 8'hc6;
assign _c_characterGenerator8x16[2282] = 8'hc6;
assign _c_characterGenerator8x16[2283] = 8'hc6;
assign _c_characterGenerator8x16[2284] = 8'h00;
assign _c_characterGenerator8x16[2285] = 8'h00;
assign _c_characterGenerator8x16[2286] = 8'h00;
assign _c_characterGenerator8x16[2287] = 8'h00;
assign _c_characterGenerator8x16[2288] = 8'h38;
assign _c_characterGenerator8x16[2289] = 8'h6c;
assign _c_characterGenerator8x16[2290] = 8'h38;
assign _c_characterGenerator8x16[2291] = 8'h00;
assign _c_characterGenerator8x16[2292] = 8'h38;
assign _c_characterGenerator8x16[2293] = 8'h6c;
assign _c_characterGenerator8x16[2294] = 8'hc6;
assign _c_characterGenerator8x16[2295] = 8'hc6;
assign _c_characterGenerator8x16[2296] = 8'hfe;
assign _c_characterGenerator8x16[2297] = 8'hc6;
assign _c_characterGenerator8x16[2298] = 8'hc6;
assign _c_characterGenerator8x16[2299] = 8'hc6;
assign _c_characterGenerator8x16[2300] = 8'h00;
assign _c_characterGenerator8x16[2301] = 8'h00;
assign _c_characterGenerator8x16[2302] = 8'h00;
assign _c_characterGenerator8x16[2303] = 8'h00;
assign _c_characterGenerator8x16[2304] = 8'h18;
assign _c_characterGenerator8x16[2305] = 8'h30;
assign _c_characterGenerator8x16[2306] = 8'h60;
assign _c_characterGenerator8x16[2307] = 8'h00;
assign _c_characterGenerator8x16[2308] = 8'hfe;
assign _c_characterGenerator8x16[2309] = 8'h66;
assign _c_characterGenerator8x16[2310] = 8'h60;
assign _c_characterGenerator8x16[2311] = 8'h7c;
assign _c_characterGenerator8x16[2312] = 8'h60;
assign _c_characterGenerator8x16[2313] = 8'h60;
assign _c_characterGenerator8x16[2314] = 8'h66;
assign _c_characterGenerator8x16[2315] = 8'hfe;
assign _c_characterGenerator8x16[2316] = 8'h00;
assign _c_characterGenerator8x16[2317] = 8'h00;
assign _c_characterGenerator8x16[2318] = 8'h00;
assign _c_characterGenerator8x16[2319] = 8'h00;
assign _c_characterGenerator8x16[2320] = 8'h00;
assign _c_characterGenerator8x16[2321] = 8'h00;
assign _c_characterGenerator8x16[2322] = 8'h00;
assign _c_characterGenerator8x16[2323] = 8'h00;
assign _c_characterGenerator8x16[2324] = 8'h00;
assign _c_characterGenerator8x16[2325] = 8'hcc;
assign _c_characterGenerator8x16[2326] = 8'h76;
assign _c_characterGenerator8x16[2327] = 8'h36;
assign _c_characterGenerator8x16[2328] = 8'h7e;
assign _c_characterGenerator8x16[2329] = 8'hd8;
assign _c_characterGenerator8x16[2330] = 8'hd8;
assign _c_characterGenerator8x16[2331] = 8'h6e;
assign _c_characterGenerator8x16[2332] = 8'h00;
assign _c_characterGenerator8x16[2333] = 8'h00;
assign _c_characterGenerator8x16[2334] = 8'h00;
assign _c_characterGenerator8x16[2335] = 8'h00;
assign _c_characterGenerator8x16[2336] = 8'h00;
assign _c_characterGenerator8x16[2337] = 8'h00;
assign _c_characterGenerator8x16[2338] = 8'h3e;
assign _c_characterGenerator8x16[2339] = 8'h6c;
assign _c_characterGenerator8x16[2340] = 8'hcc;
assign _c_characterGenerator8x16[2341] = 8'hcc;
assign _c_characterGenerator8x16[2342] = 8'hfe;
assign _c_characterGenerator8x16[2343] = 8'hcc;
assign _c_characterGenerator8x16[2344] = 8'hcc;
assign _c_characterGenerator8x16[2345] = 8'hcc;
assign _c_characterGenerator8x16[2346] = 8'hcc;
assign _c_characterGenerator8x16[2347] = 8'hce;
assign _c_characterGenerator8x16[2348] = 8'h00;
assign _c_characterGenerator8x16[2349] = 8'h00;
assign _c_characterGenerator8x16[2350] = 8'h00;
assign _c_characterGenerator8x16[2351] = 8'h00;
assign _c_characterGenerator8x16[2352] = 8'h00;
assign _c_characterGenerator8x16[2353] = 8'h10;
assign _c_characterGenerator8x16[2354] = 8'h38;
assign _c_characterGenerator8x16[2355] = 8'h6c;
assign _c_characterGenerator8x16[2356] = 8'h00;
assign _c_characterGenerator8x16[2357] = 8'h7c;
assign _c_characterGenerator8x16[2358] = 8'hc6;
assign _c_characterGenerator8x16[2359] = 8'hc6;
assign _c_characterGenerator8x16[2360] = 8'hc6;
assign _c_characterGenerator8x16[2361] = 8'hc6;
assign _c_characterGenerator8x16[2362] = 8'hc6;
assign _c_characterGenerator8x16[2363] = 8'h7c;
assign _c_characterGenerator8x16[2364] = 8'h00;
assign _c_characterGenerator8x16[2365] = 8'h00;
assign _c_characterGenerator8x16[2366] = 8'h00;
assign _c_characterGenerator8x16[2367] = 8'h00;
assign _c_characterGenerator8x16[2368] = 8'h00;
assign _c_characterGenerator8x16[2369] = 8'h00;
assign _c_characterGenerator8x16[2370] = 8'hc6;
assign _c_characterGenerator8x16[2371] = 8'h00;
assign _c_characterGenerator8x16[2372] = 8'h00;
assign _c_characterGenerator8x16[2373] = 8'h7c;
assign _c_characterGenerator8x16[2374] = 8'hc6;
assign _c_characterGenerator8x16[2375] = 8'hc6;
assign _c_characterGenerator8x16[2376] = 8'hc6;
assign _c_characterGenerator8x16[2377] = 8'hc6;
assign _c_characterGenerator8x16[2378] = 8'hc6;
assign _c_characterGenerator8x16[2379] = 8'h7c;
assign _c_characterGenerator8x16[2380] = 8'h00;
assign _c_characterGenerator8x16[2381] = 8'h00;
assign _c_characterGenerator8x16[2382] = 8'h00;
assign _c_characterGenerator8x16[2383] = 8'h00;
assign _c_characterGenerator8x16[2384] = 8'h00;
assign _c_characterGenerator8x16[2385] = 8'h60;
assign _c_characterGenerator8x16[2386] = 8'h30;
assign _c_characterGenerator8x16[2387] = 8'h18;
assign _c_characterGenerator8x16[2388] = 8'h00;
assign _c_characterGenerator8x16[2389] = 8'h7c;
assign _c_characterGenerator8x16[2390] = 8'hc6;
assign _c_characterGenerator8x16[2391] = 8'hc6;
assign _c_characterGenerator8x16[2392] = 8'hc6;
assign _c_characterGenerator8x16[2393] = 8'hc6;
assign _c_characterGenerator8x16[2394] = 8'hc6;
assign _c_characterGenerator8x16[2395] = 8'h7c;
assign _c_characterGenerator8x16[2396] = 8'h00;
assign _c_characterGenerator8x16[2397] = 8'h00;
assign _c_characterGenerator8x16[2398] = 8'h00;
assign _c_characterGenerator8x16[2399] = 8'h00;
assign _c_characterGenerator8x16[2400] = 8'h00;
assign _c_characterGenerator8x16[2401] = 8'h30;
assign _c_characterGenerator8x16[2402] = 8'h78;
assign _c_characterGenerator8x16[2403] = 8'hcc;
assign _c_characterGenerator8x16[2404] = 8'h00;
assign _c_characterGenerator8x16[2405] = 8'hcc;
assign _c_characterGenerator8x16[2406] = 8'hcc;
assign _c_characterGenerator8x16[2407] = 8'hcc;
assign _c_characterGenerator8x16[2408] = 8'hcc;
assign _c_characterGenerator8x16[2409] = 8'hcc;
assign _c_characterGenerator8x16[2410] = 8'hcc;
assign _c_characterGenerator8x16[2411] = 8'h76;
assign _c_characterGenerator8x16[2412] = 8'h00;
assign _c_characterGenerator8x16[2413] = 8'h00;
assign _c_characterGenerator8x16[2414] = 8'h00;
assign _c_characterGenerator8x16[2415] = 8'h00;
assign _c_characterGenerator8x16[2416] = 8'h00;
assign _c_characterGenerator8x16[2417] = 8'h60;
assign _c_characterGenerator8x16[2418] = 8'h30;
assign _c_characterGenerator8x16[2419] = 8'h18;
assign _c_characterGenerator8x16[2420] = 8'h00;
assign _c_characterGenerator8x16[2421] = 8'hcc;
assign _c_characterGenerator8x16[2422] = 8'hcc;
assign _c_characterGenerator8x16[2423] = 8'hcc;
assign _c_characterGenerator8x16[2424] = 8'hcc;
assign _c_characterGenerator8x16[2425] = 8'hcc;
assign _c_characterGenerator8x16[2426] = 8'hcc;
assign _c_characterGenerator8x16[2427] = 8'h76;
assign _c_characterGenerator8x16[2428] = 8'h00;
assign _c_characterGenerator8x16[2429] = 8'h00;
assign _c_characterGenerator8x16[2430] = 8'h00;
assign _c_characterGenerator8x16[2431] = 8'h00;
assign _c_characterGenerator8x16[2432] = 8'h00;
assign _c_characterGenerator8x16[2433] = 8'h00;
assign _c_characterGenerator8x16[2434] = 8'hc6;
assign _c_characterGenerator8x16[2435] = 8'h00;
assign _c_characterGenerator8x16[2436] = 8'h00;
assign _c_characterGenerator8x16[2437] = 8'hc6;
assign _c_characterGenerator8x16[2438] = 8'hc6;
assign _c_characterGenerator8x16[2439] = 8'hc6;
assign _c_characterGenerator8x16[2440] = 8'hc6;
assign _c_characterGenerator8x16[2441] = 8'hc6;
assign _c_characterGenerator8x16[2442] = 8'hc6;
assign _c_characterGenerator8x16[2443] = 8'h7e;
assign _c_characterGenerator8x16[2444] = 8'h06;
assign _c_characterGenerator8x16[2445] = 8'h0c;
assign _c_characterGenerator8x16[2446] = 8'h78;
assign _c_characterGenerator8x16[2447] = 8'h00;
assign _c_characterGenerator8x16[2448] = 8'h00;
assign _c_characterGenerator8x16[2449] = 8'hc6;
assign _c_characterGenerator8x16[2450] = 8'h00;
assign _c_characterGenerator8x16[2451] = 8'h7c;
assign _c_characterGenerator8x16[2452] = 8'hc6;
assign _c_characterGenerator8x16[2453] = 8'hc6;
assign _c_characterGenerator8x16[2454] = 8'hc6;
assign _c_characterGenerator8x16[2455] = 8'hc6;
assign _c_characterGenerator8x16[2456] = 8'hc6;
assign _c_characterGenerator8x16[2457] = 8'hc6;
assign _c_characterGenerator8x16[2458] = 8'hc6;
assign _c_characterGenerator8x16[2459] = 8'h7c;
assign _c_characterGenerator8x16[2460] = 8'h00;
assign _c_characterGenerator8x16[2461] = 8'h00;
assign _c_characterGenerator8x16[2462] = 8'h00;
assign _c_characterGenerator8x16[2463] = 8'h00;
assign _c_characterGenerator8x16[2464] = 8'h00;
assign _c_characterGenerator8x16[2465] = 8'hc6;
assign _c_characterGenerator8x16[2466] = 8'h00;
assign _c_characterGenerator8x16[2467] = 8'hc6;
assign _c_characterGenerator8x16[2468] = 8'hc6;
assign _c_characterGenerator8x16[2469] = 8'hc6;
assign _c_characterGenerator8x16[2470] = 8'hc6;
assign _c_characterGenerator8x16[2471] = 8'hc6;
assign _c_characterGenerator8x16[2472] = 8'hc6;
assign _c_characterGenerator8x16[2473] = 8'hc6;
assign _c_characterGenerator8x16[2474] = 8'hc6;
assign _c_characterGenerator8x16[2475] = 8'h7c;
assign _c_characterGenerator8x16[2476] = 8'h00;
assign _c_characterGenerator8x16[2477] = 8'h00;
assign _c_characterGenerator8x16[2478] = 8'h00;
assign _c_characterGenerator8x16[2479] = 8'h00;
assign _c_characterGenerator8x16[2480] = 8'h00;
assign _c_characterGenerator8x16[2481] = 8'h18;
assign _c_characterGenerator8x16[2482] = 8'h18;
assign _c_characterGenerator8x16[2483] = 8'h3c;
assign _c_characterGenerator8x16[2484] = 8'h66;
assign _c_characterGenerator8x16[2485] = 8'h60;
assign _c_characterGenerator8x16[2486] = 8'h60;
assign _c_characterGenerator8x16[2487] = 8'h60;
assign _c_characterGenerator8x16[2488] = 8'h66;
assign _c_characterGenerator8x16[2489] = 8'h3c;
assign _c_characterGenerator8x16[2490] = 8'h18;
assign _c_characterGenerator8x16[2491] = 8'h18;
assign _c_characterGenerator8x16[2492] = 8'h00;
assign _c_characterGenerator8x16[2493] = 8'h00;
assign _c_characterGenerator8x16[2494] = 8'h00;
assign _c_characterGenerator8x16[2495] = 8'h00;
assign _c_characterGenerator8x16[2496] = 8'h00;
assign _c_characterGenerator8x16[2497] = 8'h38;
assign _c_characterGenerator8x16[2498] = 8'h6c;
assign _c_characterGenerator8x16[2499] = 8'h64;
assign _c_characterGenerator8x16[2500] = 8'h60;
assign _c_characterGenerator8x16[2501] = 8'hf0;
assign _c_characterGenerator8x16[2502] = 8'h60;
assign _c_characterGenerator8x16[2503] = 8'h60;
assign _c_characterGenerator8x16[2504] = 8'h60;
assign _c_characterGenerator8x16[2505] = 8'h60;
assign _c_characterGenerator8x16[2506] = 8'he6;
assign _c_characterGenerator8x16[2507] = 8'hfc;
assign _c_characterGenerator8x16[2508] = 8'h00;
assign _c_characterGenerator8x16[2509] = 8'h00;
assign _c_characterGenerator8x16[2510] = 8'h00;
assign _c_characterGenerator8x16[2511] = 8'h00;
assign _c_characterGenerator8x16[2512] = 8'h00;
assign _c_characterGenerator8x16[2513] = 8'h00;
assign _c_characterGenerator8x16[2514] = 8'h66;
assign _c_characterGenerator8x16[2515] = 8'h66;
assign _c_characterGenerator8x16[2516] = 8'h3c;
assign _c_characterGenerator8x16[2517] = 8'h18;
assign _c_characterGenerator8x16[2518] = 8'h7e;
assign _c_characterGenerator8x16[2519] = 8'h18;
assign _c_characterGenerator8x16[2520] = 8'h7e;
assign _c_characterGenerator8x16[2521] = 8'h18;
assign _c_characterGenerator8x16[2522] = 8'h18;
assign _c_characterGenerator8x16[2523] = 8'h18;
assign _c_characterGenerator8x16[2524] = 8'h00;
assign _c_characterGenerator8x16[2525] = 8'h00;
assign _c_characterGenerator8x16[2526] = 8'h00;
assign _c_characterGenerator8x16[2527] = 8'h00;
assign _c_characterGenerator8x16[2528] = 8'h00;
assign _c_characterGenerator8x16[2529] = 8'hf8;
assign _c_characterGenerator8x16[2530] = 8'hcc;
assign _c_characterGenerator8x16[2531] = 8'hcc;
assign _c_characterGenerator8x16[2532] = 8'hf8;
assign _c_characterGenerator8x16[2533] = 8'hc4;
assign _c_characterGenerator8x16[2534] = 8'hcc;
assign _c_characterGenerator8x16[2535] = 8'hde;
assign _c_characterGenerator8x16[2536] = 8'hcc;
assign _c_characterGenerator8x16[2537] = 8'hcc;
assign _c_characterGenerator8x16[2538] = 8'hcc;
assign _c_characterGenerator8x16[2539] = 8'hc6;
assign _c_characterGenerator8x16[2540] = 8'h00;
assign _c_characterGenerator8x16[2541] = 8'h00;
assign _c_characterGenerator8x16[2542] = 8'h00;
assign _c_characterGenerator8x16[2543] = 8'h00;
assign _c_characterGenerator8x16[2544] = 8'h00;
assign _c_characterGenerator8x16[2545] = 8'h0e;
assign _c_characterGenerator8x16[2546] = 8'h1b;
assign _c_characterGenerator8x16[2547] = 8'h18;
assign _c_characterGenerator8x16[2548] = 8'h18;
assign _c_characterGenerator8x16[2549] = 8'h18;
assign _c_characterGenerator8x16[2550] = 8'h7e;
assign _c_characterGenerator8x16[2551] = 8'h18;
assign _c_characterGenerator8x16[2552] = 8'h18;
assign _c_characterGenerator8x16[2553] = 8'h18;
assign _c_characterGenerator8x16[2554] = 8'h18;
assign _c_characterGenerator8x16[2555] = 8'h18;
assign _c_characterGenerator8x16[2556] = 8'hd8;
assign _c_characterGenerator8x16[2557] = 8'h70;
assign _c_characterGenerator8x16[2558] = 8'h00;
assign _c_characterGenerator8x16[2559] = 8'h00;
assign _c_characterGenerator8x16[2560] = 8'h00;
assign _c_characterGenerator8x16[2561] = 8'h18;
assign _c_characterGenerator8x16[2562] = 8'h30;
assign _c_characterGenerator8x16[2563] = 8'h60;
assign _c_characterGenerator8x16[2564] = 8'h00;
assign _c_characterGenerator8x16[2565] = 8'h78;
assign _c_characterGenerator8x16[2566] = 8'h0c;
assign _c_characterGenerator8x16[2567] = 8'h7c;
assign _c_characterGenerator8x16[2568] = 8'hcc;
assign _c_characterGenerator8x16[2569] = 8'hcc;
assign _c_characterGenerator8x16[2570] = 8'hcc;
assign _c_characterGenerator8x16[2571] = 8'h76;
assign _c_characterGenerator8x16[2572] = 8'h00;
assign _c_characterGenerator8x16[2573] = 8'h00;
assign _c_characterGenerator8x16[2574] = 8'h00;
assign _c_characterGenerator8x16[2575] = 8'h00;
assign _c_characterGenerator8x16[2576] = 8'h00;
assign _c_characterGenerator8x16[2577] = 8'h0c;
assign _c_characterGenerator8x16[2578] = 8'h18;
assign _c_characterGenerator8x16[2579] = 8'h30;
assign _c_characterGenerator8x16[2580] = 8'h00;
assign _c_characterGenerator8x16[2581] = 8'h38;
assign _c_characterGenerator8x16[2582] = 8'h18;
assign _c_characterGenerator8x16[2583] = 8'h18;
assign _c_characterGenerator8x16[2584] = 8'h18;
assign _c_characterGenerator8x16[2585] = 8'h18;
assign _c_characterGenerator8x16[2586] = 8'h18;
assign _c_characterGenerator8x16[2587] = 8'h3c;
assign _c_characterGenerator8x16[2588] = 8'h00;
assign _c_characterGenerator8x16[2589] = 8'h00;
assign _c_characterGenerator8x16[2590] = 8'h00;
assign _c_characterGenerator8x16[2591] = 8'h00;
assign _c_characterGenerator8x16[2592] = 8'h00;
assign _c_characterGenerator8x16[2593] = 8'h18;
assign _c_characterGenerator8x16[2594] = 8'h30;
assign _c_characterGenerator8x16[2595] = 8'h60;
assign _c_characterGenerator8x16[2596] = 8'h00;
assign _c_characterGenerator8x16[2597] = 8'h7c;
assign _c_characterGenerator8x16[2598] = 8'hc6;
assign _c_characterGenerator8x16[2599] = 8'hc6;
assign _c_characterGenerator8x16[2600] = 8'hc6;
assign _c_characterGenerator8x16[2601] = 8'hc6;
assign _c_characterGenerator8x16[2602] = 8'hc6;
assign _c_characterGenerator8x16[2603] = 8'h7c;
assign _c_characterGenerator8x16[2604] = 8'h00;
assign _c_characterGenerator8x16[2605] = 8'h00;
assign _c_characterGenerator8x16[2606] = 8'h00;
assign _c_characterGenerator8x16[2607] = 8'h00;
assign _c_characterGenerator8x16[2608] = 8'h00;
assign _c_characterGenerator8x16[2609] = 8'h18;
assign _c_characterGenerator8x16[2610] = 8'h30;
assign _c_characterGenerator8x16[2611] = 8'h60;
assign _c_characterGenerator8x16[2612] = 8'h00;
assign _c_characterGenerator8x16[2613] = 8'hcc;
assign _c_characterGenerator8x16[2614] = 8'hcc;
assign _c_characterGenerator8x16[2615] = 8'hcc;
assign _c_characterGenerator8x16[2616] = 8'hcc;
assign _c_characterGenerator8x16[2617] = 8'hcc;
assign _c_characterGenerator8x16[2618] = 8'hcc;
assign _c_characterGenerator8x16[2619] = 8'h76;
assign _c_characterGenerator8x16[2620] = 8'h00;
assign _c_characterGenerator8x16[2621] = 8'h00;
assign _c_characterGenerator8x16[2622] = 8'h00;
assign _c_characterGenerator8x16[2623] = 8'h00;
assign _c_characterGenerator8x16[2624] = 8'h00;
assign _c_characterGenerator8x16[2625] = 8'h00;
assign _c_characterGenerator8x16[2626] = 8'h76;
assign _c_characterGenerator8x16[2627] = 8'hdc;
assign _c_characterGenerator8x16[2628] = 8'h00;
assign _c_characterGenerator8x16[2629] = 8'hdc;
assign _c_characterGenerator8x16[2630] = 8'h66;
assign _c_characterGenerator8x16[2631] = 8'h66;
assign _c_characterGenerator8x16[2632] = 8'h66;
assign _c_characterGenerator8x16[2633] = 8'h66;
assign _c_characterGenerator8x16[2634] = 8'h66;
assign _c_characterGenerator8x16[2635] = 8'h66;
assign _c_characterGenerator8x16[2636] = 8'h00;
assign _c_characterGenerator8x16[2637] = 8'h00;
assign _c_characterGenerator8x16[2638] = 8'h00;
assign _c_characterGenerator8x16[2639] = 8'h00;
assign _c_characterGenerator8x16[2640] = 8'h76;
assign _c_characterGenerator8x16[2641] = 8'hdc;
assign _c_characterGenerator8x16[2642] = 8'h00;
assign _c_characterGenerator8x16[2643] = 8'hc6;
assign _c_characterGenerator8x16[2644] = 8'he6;
assign _c_characterGenerator8x16[2645] = 8'hf6;
assign _c_characterGenerator8x16[2646] = 8'hfe;
assign _c_characterGenerator8x16[2647] = 8'hde;
assign _c_characterGenerator8x16[2648] = 8'hce;
assign _c_characterGenerator8x16[2649] = 8'hc6;
assign _c_characterGenerator8x16[2650] = 8'hc6;
assign _c_characterGenerator8x16[2651] = 8'hc6;
assign _c_characterGenerator8x16[2652] = 8'h00;
assign _c_characterGenerator8x16[2653] = 8'h00;
assign _c_characterGenerator8x16[2654] = 8'h00;
assign _c_characterGenerator8x16[2655] = 8'h00;
assign _c_characterGenerator8x16[2656] = 8'h00;
assign _c_characterGenerator8x16[2657] = 8'h3c;
assign _c_characterGenerator8x16[2658] = 8'h6c;
assign _c_characterGenerator8x16[2659] = 8'h6c;
assign _c_characterGenerator8x16[2660] = 8'h3e;
assign _c_characterGenerator8x16[2661] = 8'h00;
assign _c_characterGenerator8x16[2662] = 8'h7e;
assign _c_characterGenerator8x16[2663] = 8'h00;
assign _c_characterGenerator8x16[2664] = 8'h00;
assign _c_characterGenerator8x16[2665] = 8'h00;
assign _c_characterGenerator8x16[2666] = 8'h00;
assign _c_characterGenerator8x16[2667] = 8'h00;
assign _c_characterGenerator8x16[2668] = 8'h00;
assign _c_characterGenerator8x16[2669] = 8'h00;
assign _c_characterGenerator8x16[2670] = 8'h00;
assign _c_characterGenerator8x16[2671] = 8'h00;
assign _c_characterGenerator8x16[2672] = 8'h00;
assign _c_characterGenerator8x16[2673] = 8'h38;
assign _c_characterGenerator8x16[2674] = 8'h6c;
assign _c_characterGenerator8x16[2675] = 8'h6c;
assign _c_characterGenerator8x16[2676] = 8'h38;
assign _c_characterGenerator8x16[2677] = 8'h00;
assign _c_characterGenerator8x16[2678] = 8'h7c;
assign _c_characterGenerator8x16[2679] = 8'h00;
assign _c_characterGenerator8x16[2680] = 8'h00;
assign _c_characterGenerator8x16[2681] = 8'h00;
assign _c_characterGenerator8x16[2682] = 8'h00;
assign _c_characterGenerator8x16[2683] = 8'h00;
assign _c_characterGenerator8x16[2684] = 8'h00;
assign _c_characterGenerator8x16[2685] = 8'h00;
assign _c_characterGenerator8x16[2686] = 8'h00;
assign _c_characterGenerator8x16[2687] = 8'h00;
assign _c_characterGenerator8x16[2688] = 8'h00;
assign _c_characterGenerator8x16[2689] = 8'h00;
assign _c_characterGenerator8x16[2690] = 8'h30;
assign _c_characterGenerator8x16[2691] = 8'h30;
assign _c_characterGenerator8x16[2692] = 8'h00;
assign _c_characterGenerator8x16[2693] = 8'h30;
assign _c_characterGenerator8x16[2694] = 8'h30;
assign _c_characterGenerator8x16[2695] = 8'h60;
assign _c_characterGenerator8x16[2696] = 8'hc0;
assign _c_characterGenerator8x16[2697] = 8'hc6;
assign _c_characterGenerator8x16[2698] = 8'hc6;
assign _c_characterGenerator8x16[2699] = 8'h7c;
assign _c_characterGenerator8x16[2700] = 8'h00;
assign _c_characterGenerator8x16[2701] = 8'h00;
assign _c_characterGenerator8x16[2702] = 8'h00;
assign _c_characterGenerator8x16[2703] = 8'h00;
assign _c_characterGenerator8x16[2704] = 8'h00;
assign _c_characterGenerator8x16[2705] = 8'h00;
assign _c_characterGenerator8x16[2706] = 8'h00;
assign _c_characterGenerator8x16[2707] = 8'h00;
assign _c_characterGenerator8x16[2708] = 8'h00;
assign _c_characterGenerator8x16[2709] = 8'h00;
assign _c_characterGenerator8x16[2710] = 8'hfe;
assign _c_characterGenerator8x16[2711] = 8'hc0;
assign _c_characterGenerator8x16[2712] = 8'hc0;
assign _c_characterGenerator8x16[2713] = 8'hc0;
assign _c_characterGenerator8x16[2714] = 8'hc0;
assign _c_characterGenerator8x16[2715] = 8'h00;
assign _c_characterGenerator8x16[2716] = 8'h00;
assign _c_characterGenerator8x16[2717] = 8'h00;
assign _c_characterGenerator8x16[2718] = 8'h00;
assign _c_characterGenerator8x16[2719] = 8'h00;
assign _c_characterGenerator8x16[2720] = 8'h00;
assign _c_characterGenerator8x16[2721] = 8'h00;
assign _c_characterGenerator8x16[2722] = 8'h00;
assign _c_characterGenerator8x16[2723] = 8'h00;
assign _c_characterGenerator8x16[2724] = 8'h00;
assign _c_characterGenerator8x16[2725] = 8'h00;
assign _c_characterGenerator8x16[2726] = 8'hfe;
assign _c_characterGenerator8x16[2727] = 8'h06;
assign _c_characterGenerator8x16[2728] = 8'h06;
assign _c_characterGenerator8x16[2729] = 8'h06;
assign _c_characterGenerator8x16[2730] = 8'h06;
assign _c_characterGenerator8x16[2731] = 8'h00;
assign _c_characterGenerator8x16[2732] = 8'h00;
assign _c_characterGenerator8x16[2733] = 8'h00;
assign _c_characterGenerator8x16[2734] = 8'h00;
assign _c_characterGenerator8x16[2735] = 8'h00;
assign _c_characterGenerator8x16[2736] = 8'h00;
assign _c_characterGenerator8x16[2737] = 8'hc0;
assign _c_characterGenerator8x16[2738] = 8'hc0;
assign _c_characterGenerator8x16[2739] = 8'hc2;
assign _c_characterGenerator8x16[2740] = 8'hc6;
assign _c_characterGenerator8x16[2741] = 8'hcc;
assign _c_characterGenerator8x16[2742] = 8'h18;
assign _c_characterGenerator8x16[2743] = 8'h30;
assign _c_characterGenerator8x16[2744] = 8'h60;
assign _c_characterGenerator8x16[2745] = 8'hdc;
assign _c_characterGenerator8x16[2746] = 8'h86;
assign _c_characterGenerator8x16[2747] = 8'h0c;
assign _c_characterGenerator8x16[2748] = 8'h18;
assign _c_characterGenerator8x16[2749] = 8'h3e;
assign _c_characterGenerator8x16[2750] = 8'h00;
assign _c_characterGenerator8x16[2751] = 8'h00;
assign _c_characterGenerator8x16[2752] = 8'h00;
assign _c_characterGenerator8x16[2753] = 8'hc0;
assign _c_characterGenerator8x16[2754] = 8'hc0;
assign _c_characterGenerator8x16[2755] = 8'hc2;
assign _c_characterGenerator8x16[2756] = 8'hc6;
assign _c_characterGenerator8x16[2757] = 8'hcc;
assign _c_characterGenerator8x16[2758] = 8'h18;
assign _c_characterGenerator8x16[2759] = 8'h30;
assign _c_characterGenerator8x16[2760] = 8'h66;
assign _c_characterGenerator8x16[2761] = 8'hce;
assign _c_characterGenerator8x16[2762] = 8'h9e;
assign _c_characterGenerator8x16[2763] = 8'h3e;
assign _c_characterGenerator8x16[2764] = 8'h06;
assign _c_characterGenerator8x16[2765] = 8'h06;
assign _c_characterGenerator8x16[2766] = 8'h00;
assign _c_characterGenerator8x16[2767] = 8'h00;
assign _c_characterGenerator8x16[2768] = 8'h00;
assign _c_characterGenerator8x16[2769] = 8'h00;
assign _c_characterGenerator8x16[2770] = 8'h18;
assign _c_characterGenerator8x16[2771] = 8'h18;
assign _c_characterGenerator8x16[2772] = 8'h00;
assign _c_characterGenerator8x16[2773] = 8'h18;
assign _c_characterGenerator8x16[2774] = 8'h18;
assign _c_characterGenerator8x16[2775] = 8'h18;
assign _c_characterGenerator8x16[2776] = 8'h3c;
assign _c_characterGenerator8x16[2777] = 8'h3c;
assign _c_characterGenerator8x16[2778] = 8'h3c;
assign _c_characterGenerator8x16[2779] = 8'h18;
assign _c_characterGenerator8x16[2780] = 8'h00;
assign _c_characterGenerator8x16[2781] = 8'h00;
assign _c_characterGenerator8x16[2782] = 8'h00;
assign _c_characterGenerator8x16[2783] = 8'h00;
assign _c_characterGenerator8x16[2784] = 8'h00;
assign _c_characterGenerator8x16[2785] = 8'h00;
assign _c_characterGenerator8x16[2786] = 8'h00;
assign _c_characterGenerator8x16[2787] = 8'h00;
assign _c_characterGenerator8x16[2788] = 8'h00;
assign _c_characterGenerator8x16[2789] = 8'h36;
assign _c_characterGenerator8x16[2790] = 8'h6c;
assign _c_characterGenerator8x16[2791] = 8'hd8;
assign _c_characterGenerator8x16[2792] = 8'h6c;
assign _c_characterGenerator8x16[2793] = 8'h36;
assign _c_characterGenerator8x16[2794] = 8'h00;
assign _c_characterGenerator8x16[2795] = 8'h00;
assign _c_characterGenerator8x16[2796] = 8'h00;
assign _c_characterGenerator8x16[2797] = 8'h00;
assign _c_characterGenerator8x16[2798] = 8'h00;
assign _c_characterGenerator8x16[2799] = 8'h00;
assign _c_characterGenerator8x16[2800] = 8'h00;
assign _c_characterGenerator8x16[2801] = 8'h00;
assign _c_characterGenerator8x16[2802] = 8'h00;
assign _c_characterGenerator8x16[2803] = 8'h00;
assign _c_characterGenerator8x16[2804] = 8'h00;
assign _c_characterGenerator8x16[2805] = 8'hd8;
assign _c_characterGenerator8x16[2806] = 8'h6c;
assign _c_characterGenerator8x16[2807] = 8'h36;
assign _c_characterGenerator8x16[2808] = 8'h6c;
assign _c_characterGenerator8x16[2809] = 8'hd8;
assign _c_characterGenerator8x16[2810] = 8'h00;
assign _c_characterGenerator8x16[2811] = 8'h00;
assign _c_characterGenerator8x16[2812] = 8'h00;
assign _c_characterGenerator8x16[2813] = 8'h00;
assign _c_characterGenerator8x16[2814] = 8'h00;
assign _c_characterGenerator8x16[2815] = 8'h00;
assign _c_characterGenerator8x16[2816] = 8'h11;
assign _c_characterGenerator8x16[2817] = 8'h44;
assign _c_characterGenerator8x16[2818] = 8'h11;
assign _c_characterGenerator8x16[2819] = 8'h44;
assign _c_characterGenerator8x16[2820] = 8'h11;
assign _c_characterGenerator8x16[2821] = 8'h44;
assign _c_characterGenerator8x16[2822] = 8'h11;
assign _c_characterGenerator8x16[2823] = 8'h44;
assign _c_characterGenerator8x16[2824] = 8'h11;
assign _c_characterGenerator8x16[2825] = 8'h44;
assign _c_characterGenerator8x16[2826] = 8'h11;
assign _c_characterGenerator8x16[2827] = 8'h44;
assign _c_characterGenerator8x16[2828] = 8'h11;
assign _c_characterGenerator8x16[2829] = 8'h44;
assign _c_characterGenerator8x16[2830] = 8'h11;
assign _c_characterGenerator8x16[2831] = 8'h44;
assign _c_characterGenerator8x16[2832] = 8'h55;
assign _c_characterGenerator8x16[2833] = 8'haa;
assign _c_characterGenerator8x16[2834] = 8'h55;
assign _c_characterGenerator8x16[2835] = 8'haa;
assign _c_characterGenerator8x16[2836] = 8'h55;
assign _c_characterGenerator8x16[2837] = 8'haa;
assign _c_characterGenerator8x16[2838] = 8'h55;
assign _c_characterGenerator8x16[2839] = 8'haa;
assign _c_characterGenerator8x16[2840] = 8'h55;
assign _c_characterGenerator8x16[2841] = 8'haa;
assign _c_characterGenerator8x16[2842] = 8'h55;
assign _c_characterGenerator8x16[2843] = 8'haa;
assign _c_characterGenerator8x16[2844] = 8'h55;
assign _c_characterGenerator8x16[2845] = 8'haa;
assign _c_characterGenerator8x16[2846] = 8'h55;
assign _c_characterGenerator8x16[2847] = 8'haa;
assign _c_characterGenerator8x16[2848] = 8'hdd;
assign _c_characterGenerator8x16[2849] = 8'h77;
assign _c_characterGenerator8x16[2850] = 8'hdd;
assign _c_characterGenerator8x16[2851] = 8'h77;
assign _c_characterGenerator8x16[2852] = 8'hdd;
assign _c_characterGenerator8x16[2853] = 8'h77;
assign _c_characterGenerator8x16[2854] = 8'hdd;
assign _c_characterGenerator8x16[2855] = 8'h77;
assign _c_characterGenerator8x16[2856] = 8'hdd;
assign _c_characterGenerator8x16[2857] = 8'h77;
assign _c_characterGenerator8x16[2858] = 8'hdd;
assign _c_characterGenerator8x16[2859] = 8'h77;
assign _c_characterGenerator8x16[2860] = 8'hdd;
assign _c_characterGenerator8x16[2861] = 8'h77;
assign _c_characterGenerator8x16[2862] = 8'hdd;
assign _c_characterGenerator8x16[2863] = 8'h77;
assign _c_characterGenerator8x16[2864] = 8'h18;
assign _c_characterGenerator8x16[2865] = 8'h18;
assign _c_characterGenerator8x16[2866] = 8'h18;
assign _c_characterGenerator8x16[2867] = 8'h18;
assign _c_characterGenerator8x16[2868] = 8'h18;
assign _c_characterGenerator8x16[2869] = 8'h18;
assign _c_characterGenerator8x16[2870] = 8'h18;
assign _c_characterGenerator8x16[2871] = 8'h18;
assign _c_characterGenerator8x16[2872] = 8'h18;
assign _c_characterGenerator8x16[2873] = 8'h18;
assign _c_characterGenerator8x16[2874] = 8'h18;
assign _c_characterGenerator8x16[2875] = 8'h18;
assign _c_characterGenerator8x16[2876] = 8'h18;
assign _c_characterGenerator8x16[2877] = 8'h18;
assign _c_characterGenerator8x16[2878] = 8'h18;
assign _c_characterGenerator8x16[2879] = 8'h18;
assign _c_characterGenerator8x16[2880] = 8'h18;
assign _c_characterGenerator8x16[2881] = 8'h18;
assign _c_characterGenerator8x16[2882] = 8'h18;
assign _c_characterGenerator8x16[2883] = 8'h18;
assign _c_characterGenerator8x16[2884] = 8'h18;
assign _c_characterGenerator8x16[2885] = 8'h18;
assign _c_characterGenerator8x16[2886] = 8'h18;
assign _c_characterGenerator8x16[2887] = 8'hf8;
assign _c_characterGenerator8x16[2888] = 8'h18;
assign _c_characterGenerator8x16[2889] = 8'h18;
assign _c_characterGenerator8x16[2890] = 8'h18;
assign _c_characterGenerator8x16[2891] = 8'h18;
assign _c_characterGenerator8x16[2892] = 8'h18;
assign _c_characterGenerator8x16[2893] = 8'h18;
assign _c_characterGenerator8x16[2894] = 8'h18;
assign _c_characterGenerator8x16[2895] = 8'h18;
assign _c_characterGenerator8x16[2896] = 8'h18;
assign _c_characterGenerator8x16[2897] = 8'h18;
assign _c_characterGenerator8x16[2898] = 8'h18;
assign _c_characterGenerator8x16[2899] = 8'h18;
assign _c_characterGenerator8x16[2900] = 8'h18;
assign _c_characterGenerator8x16[2901] = 8'hf8;
assign _c_characterGenerator8x16[2902] = 8'h18;
assign _c_characterGenerator8x16[2903] = 8'hf8;
assign _c_characterGenerator8x16[2904] = 8'h18;
assign _c_characterGenerator8x16[2905] = 8'h18;
assign _c_characterGenerator8x16[2906] = 8'h18;
assign _c_characterGenerator8x16[2907] = 8'h18;
assign _c_characterGenerator8x16[2908] = 8'h18;
assign _c_characterGenerator8x16[2909] = 8'h18;
assign _c_characterGenerator8x16[2910] = 8'h18;
assign _c_characterGenerator8x16[2911] = 8'h18;
assign _c_characterGenerator8x16[2912] = 8'h36;
assign _c_characterGenerator8x16[2913] = 8'h36;
assign _c_characterGenerator8x16[2914] = 8'h36;
assign _c_characterGenerator8x16[2915] = 8'h36;
assign _c_characterGenerator8x16[2916] = 8'h36;
assign _c_characterGenerator8x16[2917] = 8'h36;
assign _c_characterGenerator8x16[2918] = 8'h36;
assign _c_characterGenerator8x16[2919] = 8'hf6;
assign _c_characterGenerator8x16[2920] = 8'h36;
assign _c_characterGenerator8x16[2921] = 8'h36;
assign _c_characterGenerator8x16[2922] = 8'h36;
assign _c_characterGenerator8x16[2923] = 8'h36;
assign _c_characterGenerator8x16[2924] = 8'h36;
assign _c_characterGenerator8x16[2925] = 8'h36;
assign _c_characterGenerator8x16[2926] = 8'h36;
assign _c_characterGenerator8x16[2927] = 8'h36;
assign _c_characterGenerator8x16[2928] = 8'h00;
assign _c_characterGenerator8x16[2929] = 8'h00;
assign _c_characterGenerator8x16[2930] = 8'h00;
assign _c_characterGenerator8x16[2931] = 8'h00;
assign _c_characterGenerator8x16[2932] = 8'h00;
assign _c_characterGenerator8x16[2933] = 8'h00;
assign _c_characterGenerator8x16[2934] = 8'h00;
assign _c_characterGenerator8x16[2935] = 8'hfe;
assign _c_characterGenerator8x16[2936] = 8'h36;
assign _c_characterGenerator8x16[2937] = 8'h36;
assign _c_characterGenerator8x16[2938] = 8'h36;
assign _c_characterGenerator8x16[2939] = 8'h36;
assign _c_characterGenerator8x16[2940] = 8'h36;
assign _c_characterGenerator8x16[2941] = 8'h36;
assign _c_characterGenerator8x16[2942] = 8'h36;
assign _c_characterGenerator8x16[2943] = 8'h36;
assign _c_characterGenerator8x16[2944] = 8'h00;
assign _c_characterGenerator8x16[2945] = 8'h00;
assign _c_characterGenerator8x16[2946] = 8'h00;
assign _c_characterGenerator8x16[2947] = 8'h00;
assign _c_characterGenerator8x16[2948] = 8'h00;
assign _c_characterGenerator8x16[2949] = 8'hf8;
assign _c_characterGenerator8x16[2950] = 8'h18;
assign _c_characterGenerator8x16[2951] = 8'hf8;
assign _c_characterGenerator8x16[2952] = 8'h18;
assign _c_characterGenerator8x16[2953] = 8'h18;
assign _c_characterGenerator8x16[2954] = 8'h18;
assign _c_characterGenerator8x16[2955] = 8'h18;
assign _c_characterGenerator8x16[2956] = 8'h18;
assign _c_characterGenerator8x16[2957] = 8'h18;
assign _c_characterGenerator8x16[2958] = 8'h18;
assign _c_characterGenerator8x16[2959] = 8'h18;
assign _c_characterGenerator8x16[2960] = 8'h36;
assign _c_characterGenerator8x16[2961] = 8'h36;
assign _c_characterGenerator8x16[2962] = 8'h36;
assign _c_characterGenerator8x16[2963] = 8'h36;
assign _c_characterGenerator8x16[2964] = 8'h36;
assign _c_characterGenerator8x16[2965] = 8'hf6;
assign _c_characterGenerator8x16[2966] = 8'h06;
assign _c_characterGenerator8x16[2967] = 8'hf6;
assign _c_characterGenerator8x16[2968] = 8'h36;
assign _c_characterGenerator8x16[2969] = 8'h36;
assign _c_characterGenerator8x16[2970] = 8'h36;
assign _c_characterGenerator8x16[2971] = 8'h36;
assign _c_characterGenerator8x16[2972] = 8'h36;
assign _c_characterGenerator8x16[2973] = 8'h36;
assign _c_characterGenerator8x16[2974] = 8'h36;
assign _c_characterGenerator8x16[2975] = 8'h36;
assign _c_characterGenerator8x16[2976] = 8'h36;
assign _c_characterGenerator8x16[2977] = 8'h36;
assign _c_characterGenerator8x16[2978] = 8'h36;
assign _c_characterGenerator8x16[2979] = 8'h36;
assign _c_characterGenerator8x16[2980] = 8'h36;
assign _c_characterGenerator8x16[2981] = 8'h36;
assign _c_characterGenerator8x16[2982] = 8'h36;
assign _c_characterGenerator8x16[2983] = 8'h36;
assign _c_characterGenerator8x16[2984] = 8'h36;
assign _c_characterGenerator8x16[2985] = 8'h36;
assign _c_characterGenerator8x16[2986] = 8'h36;
assign _c_characterGenerator8x16[2987] = 8'h36;
assign _c_characterGenerator8x16[2988] = 8'h36;
assign _c_characterGenerator8x16[2989] = 8'h36;
assign _c_characterGenerator8x16[2990] = 8'h36;
assign _c_characterGenerator8x16[2991] = 8'h36;
assign _c_characterGenerator8x16[2992] = 8'h00;
assign _c_characterGenerator8x16[2993] = 8'h00;
assign _c_characterGenerator8x16[2994] = 8'h00;
assign _c_characterGenerator8x16[2995] = 8'h00;
assign _c_characterGenerator8x16[2996] = 8'h00;
assign _c_characterGenerator8x16[2997] = 8'hfe;
assign _c_characterGenerator8x16[2998] = 8'h06;
assign _c_characterGenerator8x16[2999] = 8'hf6;
assign _c_characterGenerator8x16[3000] = 8'h36;
assign _c_characterGenerator8x16[3001] = 8'h36;
assign _c_characterGenerator8x16[3002] = 8'h36;
assign _c_characterGenerator8x16[3003] = 8'h36;
assign _c_characterGenerator8x16[3004] = 8'h36;
assign _c_characterGenerator8x16[3005] = 8'h36;
assign _c_characterGenerator8x16[3006] = 8'h36;
assign _c_characterGenerator8x16[3007] = 8'h36;
assign _c_characterGenerator8x16[3008] = 8'h36;
assign _c_characterGenerator8x16[3009] = 8'h36;
assign _c_characterGenerator8x16[3010] = 8'h36;
assign _c_characterGenerator8x16[3011] = 8'h36;
assign _c_characterGenerator8x16[3012] = 8'h36;
assign _c_characterGenerator8x16[3013] = 8'hf6;
assign _c_characterGenerator8x16[3014] = 8'h06;
assign _c_characterGenerator8x16[3015] = 8'hfe;
assign _c_characterGenerator8x16[3016] = 8'h00;
assign _c_characterGenerator8x16[3017] = 8'h00;
assign _c_characterGenerator8x16[3018] = 8'h00;
assign _c_characterGenerator8x16[3019] = 8'h00;
assign _c_characterGenerator8x16[3020] = 8'h00;
assign _c_characterGenerator8x16[3021] = 8'h00;
assign _c_characterGenerator8x16[3022] = 8'h00;
assign _c_characterGenerator8x16[3023] = 8'h00;
assign _c_characterGenerator8x16[3024] = 8'h36;
assign _c_characterGenerator8x16[3025] = 8'h36;
assign _c_characterGenerator8x16[3026] = 8'h36;
assign _c_characterGenerator8x16[3027] = 8'h36;
assign _c_characterGenerator8x16[3028] = 8'h36;
assign _c_characterGenerator8x16[3029] = 8'h36;
assign _c_characterGenerator8x16[3030] = 8'h36;
assign _c_characterGenerator8x16[3031] = 8'hfe;
assign _c_characterGenerator8x16[3032] = 8'h00;
assign _c_characterGenerator8x16[3033] = 8'h00;
assign _c_characterGenerator8x16[3034] = 8'h00;
assign _c_characterGenerator8x16[3035] = 8'h00;
assign _c_characterGenerator8x16[3036] = 8'h00;
assign _c_characterGenerator8x16[3037] = 8'h00;
assign _c_characterGenerator8x16[3038] = 8'h00;
assign _c_characterGenerator8x16[3039] = 8'h00;
assign _c_characterGenerator8x16[3040] = 8'h18;
assign _c_characterGenerator8x16[3041] = 8'h18;
assign _c_characterGenerator8x16[3042] = 8'h18;
assign _c_characterGenerator8x16[3043] = 8'h18;
assign _c_characterGenerator8x16[3044] = 8'h18;
assign _c_characterGenerator8x16[3045] = 8'hf8;
assign _c_characterGenerator8x16[3046] = 8'h18;
assign _c_characterGenerator8x16[3047] = 8'hf8;
assign _c_characterGenerator8x16[3048] = 8'h00;
assign _c_characterGenerator8x16[3049] = 8'h00;
assign _c_characterGenerator8x16[3050] = 8'h00;
assign _c_characterGenerator8x16[3051] = 8'h00;
assign _c_characterGenerator8x16[3052] = 8'h00;
assign _c_characterGenerator8x16[3053] = 8'h00;
assign _c_characterGenerator8x16[3054] = 8'h00;
assign _c_characterGenerator8x16[3055] = 8'h00;
assign _c_characterGenerator8x16[3056] = 8'h00;
assign _c_characterGenerator8x16[3057] = 8'h00;
assign _c_characterGenerator8x16[3058] = 8'h00;
assign _c_characterGenerator8x16[3059] = 8'h00;
assign _c_characterGenerator8x16[3060] = 8'h00;
assign _c_characterGenerator8x16[3061] = 8'h00;
assign _c_characterGenerator8x16[3062] = 8'h00;
assign _c_characterGenerator8x16[3063] = 8'hf8;
assign _c_characterGenerator8x16[3064] = 8'h18;
assign _c_characterGenerator8x16[3065] = 8'h18;
assign _c_characterGenerator8x16[3066] = 8'h18;
assign _c_characterGenerator8x16[3067] = 8'h18;
assign _c_characterGenerator8x16[3068] = 8'h18;
assign _c_characterGenerator8x16[3069] = 8'h18;
assign _c_characterGenerator8x16[3070] = 8'h18;
assign _c_characterGenerator8x16[3071] = 8'h18;
assign _c_characterGenerator8x16[3072] = 8'h18;
assign _c_characterGenerator8x16[3073] = 8'h18;
assign _c_characterGenerator8x16[3074] = 8'h18;
assign _c_characterGenerator8x16[3075] = 8'h18;
assign _c_characterGenerator8x16[3076] = 8'h18;
assign _c_characterGenerator8x16[3077] = 8'h18;
assign _c_characterGenerator8x16[3078] = 8'h18;
assign _c_characterGenerator8x16[3079] = 8'h1f;
assign _c_characterGenerator8x16[3080] = 8'h00;
assign _c_characterGenerator8x16[3081] = 8'h00;
assign _c_characterGenerator8x16[3082] = 8'h00;
assign _c_characterGenerator8x16[3083] = 8'h00;
assign _c_characterGenerator8x16[3084] = 8'h00;
assign _c_characterGenerator8x16[3085] = 8'h00;
assign _c_characterGenerator8x16[3086] = 8'h00;
assign _c_characterGenerator8x16[3087] = 8'h00;
assign _c_characterGenerator8x16[3088] = 8'h18;
assign _c_characterGenerator8x16[3089] = 8'h18;
assign _c_characterGenerator8x16[3090] = 8'h18;
assign _c_characterGenerator8x16[3091] = 8'h18;
assign _c_characterGenerator8x16[3092] = 8'h18;
assign _c_characterGenerator8x16[3093] = 8'h18;
assign _c_characterGenerator8x16[3094] = 8'h18;
assign _c_characterGenerator8x16[3095] = 8'hff;
assign _c_characterGenerator8x16[3096] = 8'h00;
assign _c_characterGenerator8x16[3097] = 8'h00;
assign _c_characterGenerator8x16[3098] = 8'h00;
assign _c_characterGenerator8x16[3099] = 8'h00;
assign _c_characterGenerator8x16[3100] = 8'h00;
assign _c_characterGenerator8x16[3101] = 8'h00;
assign _c_characterGenerator8x16[3102] = 8'h00;
assign _c_characterGenerator8x16[3103] = 8'h00;
assign _c_characterGenerator8x16[3104] = 8'h00;
assign _c_characterGenerator8x16[3105] = 8'h00;
assign _c_characterGenerator8x16[3106] = 8'h00;
assign _c_characterGenerator8x16[3107] = 8'h00;
assign _c_characterGenerator8x16[3108] = 8'h00;
assign _c_characterGenerator8x16[3109] = 8'h00;
assign _c_characterGenerator8x16[3110] = 8'h00;
assign _c_characterGenerator8x16[3111] = 8'hff;
assign _c_characterGenerator8x16[3112] = 8'h18;
assign _c_characterGenerator8x16[3113] = 8'h18;
assign _c_characterGenerator8x16[3114] = 8'h18;
assign _c_characterGenerator8x16[3115] = 8'h18;
assign _c_characterGenerator8x16[3116] = 8'h18;
assign _c_characterGenerator8x16[3117] = 8'h18;
assign _c_characterGenerator8x16[3118] = 8'h18;
assign _c_characterGenerator8x16[3119] = 8'h18;
assign _c_characterGenerator8x16[3120] = 8'h18;
assign _c_characterGenerator8x16[3121] = 8'h18;
assign _c_characterGenerator8x16[3122] = 8'h18;
assign _c_characterGenerator8x16[3123] = 8'h18;
assign _c_characterGenerator8x16[3124] = 8'h18;
assign _c_characterGenerator8x16[3125] = 8'h18;
assign _c_characterGenerator8x16[3126] = 8'h18;
assign _c_characterGenerator8x16[3127] = 8'h1f;
assign _c_characterGenerator8x16[3128] = 8'h18;
assign _c_characterGenerator8x16[3129] = 8'h18;
assign _c_characterGenerator8x16[3130] = 8'h18;
assign _c_characterGenerator8x16[3131] = 8'h18;
assign _c_characterGenerator8x16[3132] = 8'h18;
assign _c_characterGenerator8x16[3133] = 8'h18;
assign _c_characterGenerator8x16[3134] = 8'h18;
assign _c_characterGenerator8x16[3135] = 8'h18;
assign _c_characterGenerator8x16[3136] = 8'h00;
assign _c_characterGenerator8x16[3137] = 8'h00;
assign _c_characterGenerator8x16[3138] = 8'h00;
assign _c_characterGenerator8x16[3139] = 8'h00;
assign _c_characterGenerator8x16[3140] = 8'h00;
assign _c_characterGenerator8x16[3141] = 8'h00;
assign _c_characterGenerator8x16[3142] = 8'h00;
assign _c_characterGenerator8x16[3143] = 8'hff;
assign _c_characterGenerator8x16[3144] = 8'h00;
assign _c_characterGenerator8x16[3145] = 8'h00;
assign _c_characterGenerator8x16[3146] = 8'h00;
assign _c_characterGenerator8x16[3147] = 8'h00;
assign _c_characterGenerator8x16[3148] = 8'h00;
assign _c_characterGenerator8x16[3149] = 8'h00;
assign _c_characterGenerator8x16[3150] = 8'h00;
assign _c_characterGenerator8x16[3151] = 8'h00;
assign _c_characterGenerator8x16[3152] = 8'h18;
assign _c_characterGenerator8x16[3153] = 8'h18;
assign _c_characterGenerator8x16[3154] = 8'h18;
assign _c_characterGenerator8x16[3155] = 8'h18;
assign _c_characterGenerator8x16[3156] = 8'h18;
assign _c_characterGenerator8x16[3157] = 8'h18;
assign _c_characterGenerator8x16[3158] = 8'h18;
assign _c_characterGenerator8x16[3159] = 8'hff;
assign _c_characterGenerator8x16[3160] = 8'h18;
assign _c_characterGenerator8x16[3161] = 8'h18;
assign _c_characterGenerator8x16[3162] = 8'h18;
assign _c_characterGenerator8x16[3163] = 8'h18;
assign _c_characterGenerator8x16[3164] = 8'h18;
assign _c_characterGenerator8x16[3165] = 8'h18;
assign _c_characterGenerator8x16[3166] = 8'h18;
assign _c_characterGenerator8x16[3167] = 8'h18;
assign _c_characterGenerator8x16[3168] = 8'h18;
assign _c_characterGenerator8x16[3169] = 8'h18;
assign _c_characterGenerator8x16[3170] = 8'h18;
assign _c_characterGenerator8x16[3171] = 8'h18;
assign _c_characterGenerator8x16[3172] = 8'h18;
assign _c_characterGenerator8x16[3173] = 8'h1f;
assign _c_characterGenerator8x16[3174] = 8'h18;
assign _c_characterGenerator8x16[3175] = 8'h1f;
assign _c_characterGenerator8x16[3176] = 8'h18;
assign _c_characterGenerator8x16[3177] = 8'h18;
assign _c_characterGenerator8x16[3178] = 8'h18;
assign _c_characterGenerator8x16[3179] = 8'h18;
assign _c_characterGenerator8x16[3180] = 8'h18;
assign _c_characterGenerator8x16[3181] = 8'h18;
assign _c_characterGenerator8x16[3182] = 8'h18;
assign _c_characterGenerator8x16[3183] = 8'h18;
assign _c_characterGenerator8x16[3184] = 8'h36;
assign _c_characterGenerator8x16[3185] = 8'h36;
assign _c_characterGenerator8x16[3186] = 8'h36;
assign _c_characterGenerator8x16[3187] = 8'h36;
assign _c_characterGenerator8x16[3188] = 8'h36;
assign _c_characterGenerator8x16[3189] = 8'h36;
assign _c_characterGenerator8x16[3190] = 8'h36;
assign _c_characterGenerator8x16[3191] = 8'h37;
assign _c_characterGenerator8x16[3192] = 8'h36;
assign _c_characterGenerator8x16[3193] = 8'h36;
assign _c_characterGenerator8x16[3194] = 8'h36;
assign _c_characterGenerator8x16[3195] = 8'h36;
assign _c_characterGenerator8x16[3196] = 8'h36;
assign _c_characterGenerator8x16[3197] = 8'h36;
assign _c_characterGenerator8x16[3198] = 8'h36;
assign _c_characterGenerator8x16[3199] = 8'h36;
assign _c_characterGenerator8x16[3200] = 8'h36;
assign _c_characterGenerator8x16[3201] = 8'h36;
assign _c_characterGenerator8x16[3202] = 8'h36;
assign _c_characterGenerator8x16[3203] = 8'h36;
assign _c_characterGenerator8x16[3204] = 8'h36;
assign _c_characterGenerator8x16[3205] = 8'h37;
assign _c_characterGenerator8x16[3206] = 8'h30;
assign _c_characterGenerator8x16[3207] = 8'h3f;
assign _c_characterGenerator8x16[3208] = 8'h00;
assign _c_characterGenerator8x16[3209] = 8'h00;
assign _c_characterGenerator8x16[3210] = 8'h00;
assign _c_characterGenerator8x16[3211] = 8'h00;
assign _c_characterGenerator8x16[3212] = 8'h00;
assign _c_characterGenerator8x16[3213] = 8'h00;
assign _c_characterGenerator8x16[3214] = 8'h00;
assign _c_characterGenerator8x16[3215] = 8'h00;
assign _c_characterGenerator8x16[3216] = 8'h00;
assign _c_characterGenerator8x16[3217] = 8'h00;
assign _c_characterGenerator8x16[3218] = 8'h00;
assign _c_characterGenerator8x16[3219] = 8'h00;
assign _c_characterGenerator8x16[3220] = 8'h00;
assign _c_characterGenerator8x16[3221] = 8'h3f;
assign _c_characterGenerator8x16[3222] = 8'h30;
assign _c_characterGenerator8x16[3223] = 8'h37;
assign _c_characterGenerator8x16[3224] = 8'h36;
assign _c_characterGenerator8x16[3225] = 8'h36;
assign _c_characterGenerator8x16[3226] = 8'h36;
assign _c_characterGenerator8x16[3227] = 8'h36;
assign _c_characterGenerator8x16[3228] = 8'h36;
assign _c_characterGenerator8x16[3229] = 8'h36;
assign _c_characterGenerator8x16[3230] = 8'h36;
assign _c_characterGenerator8x16[3231] = 8'h36;
assign _c_characterGenerator8x16[3232] = 8'h36;
assign _c_characterGenerator8x16[3233] = 8'h36;
assign _c_characterGenerator8x16[3234] = 8'h36;
assign _c_characterGenerator8x16[3235] = 8'h36;
assign _c_characterGenerator8x16[3236] = 8'h36;
assign _c_characterGenerator8x16[3237] = 8'hf7;
assign _c_characterGenerator8x16[3238] = 8'h00;
assign _c_characterGenerator8x16[3239] = 8'hff;
assign _c_characterGenerator8x16[3240] = 8'h00;
assign _c_characterGenerator8x16[3241] = 8'h00;
assign _c_characterGenerator8x16[3242] = 8'h00;
assign _c_characterGenerator8x16[3243] = 8'h00;
assign _c_characterGenerator8x16[3244] = 8'h00;
assign _c_characterGenerator8x16[3245] = 8'h00;
assign _c_characterGenerator8x16[3246] = 8'h00;
assign _c_characterGenerator8x16[3247] = 8'h00;
assign _c_characterGenerator8x16[3248] = 8'h00;
assign _c_characterGenerator8x16[3249] = 8'h00;
assign _c_characterGenerator8x16[3250] = 8'h00;
assign _c_characterGenerator8x16[3251] = 8'h00;
assign _c_characterGenerator8x16[3252] = 8'h00;
assign _c_characterGenerator8x16[3253] = 8'hff;
assign _c_characterGenerator8x16[3254] = 8'h00;
assign _c_characterGenerator8x16[3255] = 8'hf7;
assign _c_characterGenerator8x16[3256] = 8'h36;
assign _c_characterGenerator8x16[3257] = 8'h36;
assign _c_characterGenerator8x16[3258] = 8'h36;
assign _c_characterGenerator8x16[3259] = 8'h36;
assign _c_characterGenerator8x16[3260] = 8'h36;
assign _c_characterGenerator8x16[3261] = 8'h36;
assign _c_characterGenerator8x16[3262] = 8'h36;
assign _c_characterGenerator8x16[3263] = 8'h36;
assign _c_characterGenerator8x16[3264] = 8'h36;
assign _c_characterGenerator8x16[3265] = 8'h36;
assign _c_characterGenerator8x16[3266] = 8'h36;
assign _c_characterGenerator8x16[3267] = 8'h36;
assign _c_characterGenerator8x16[3268] = 8'h36;
assign _c_characterGenerator8x16[3269] = 8'h37;
assign _c_characterGenerator8x16[3270] = 8'h30;
assign _c_characterGenerator8x16[3271] = 8'h37;
assign _c_characterGenerator8x16[3272] = 8'h36;
assign _c_characterGenerator8x16[3273] = 8'h36;
assign _c_characterGenerator8x16[3274] = 8'h36;
assign _c_characterGenerator8x16[3275] = 8'h36;
assign _c_characterGenerator8x16[3276] = 8'h36;
assign _c_characterGenerator8x16[3277] = 8'h36;
assign _c_characterGenerator8x16[3278] = 8'h36;
assign _c_characterGenerator8x16[3279] = 8'h36;
assign _c_characterGenerator8x16[3280] = 8'h00;
assign _c_characterGenerator8x16[3281] = 8'h00;
assign _c_characterGenerator8x16[3282] = 8'h00;
assign _c_characterGenerator8x16[3283] = 8'h00;
assign _c_characterGenerator8x16[3284] = 8'h00;
assign _c_characterGenerator8x16[3285] = 8'hff;
assign _c_characterGenerator8x16[3286] = 8'h00;
assign _c_characterGenerator8x16[3287] = 8'hff;
assign _c_characterGenerator8x16[3288] = 8'h00;
assign _c_characterGenerator8x16[3289] = 8'h00;
assign _c_characterGenerator8x16[3290] = 8'h00;
assign _c_characterGenerator8x16[3291] = 8'h00;
assign _c_characterGenerator8x16[3292] = 8'h00;
assign _c_characterGenerator8x16[3293] = 8'h00;
assign _c_characterGenerator8x16[3294] = 8'h00;
assign _c_characterGenerator8x16[3295] = 8'h00;
assign _c_characterGenerator8x16[3296] = 8'h36;
assign _c_characterGenerator8x16[3297] = 8'h36;
assign _c_characterGenerator8x16[3298] = 8'h36;
assign _c_characterGenerator8x16[3299] = 8'h36;
assign _c_characterGenerator8x16[3300] = 8'h36;
assign _c_characterGenerator8x16[3301] = 8'hf7;
assign _c_characterGenerator8x16[3302] = 8'h00;
assign _c_characterGenerator8x16[3303] = 8'hf7;
assign _c_characterGenerator8x16[3304] = 8'h36;
assign _c_characterGenerator8x16[3305] = 8'h36;
assign _c_characterGenerator8x16[3306] = 8'h36;
assign _c_characterGenerator8x16[3307] = 8'h36;
assign _c_characterGenerator8x16[3308] = 8'h36;
assign _c_characterGenerator8x16[3309] = 8'h36;
assign _c_characterGenerator8x16[3310] = 8'h36;
assign _c_characterGenerator8x16[3311] = 8'h36;
assign _c_characterGenerator8x16[3312] = 8'h18;
assign _c_characterGenerator8x16[3313] = 8'h18;
assign _c_characterGenerator8x16[3314] = 8'h18;
assign _c_characterGenerator8x16[3315] = 8'h18;
assign _c_characterGenerator8x16[3316] = 8'h18;
assign _c_characterGenerator8x16[3317] = 8'hff;
assign _c_characterGenerator8x16[3318] = 8'h00;
assign _c_characterGenerator8x16[3319] = 8'hff;
assign _c_characterGenerator8x16[3320] = 8'h00;
assign _c_characterGenerator8x16[3321] = 8'h00;
assign _c_characterGenerator8x16[3322] = 8'h00;
assign _c_characterGenerator8x16[3323] = 8'h00;
assign _c_characterGenerator8x16[3324] = 8'h00;
assign _c_characterGenerator8x16[3325] = 8'h00;
assign _c_characterGenerator8x16[3326] = 8'h00;
assign _c_characterGenerator8x16[3327] = 8'h00;
assign _c_characterGenerator8x16[3328] = 8'h36;
assign _c_characterGenerator8x16[3329] = 8'h36;
assign _c_characterGenerator8x16[3330] = 8'h36;
assign _c_characterGenerator8x16[3331] = 8'h36;
assign _c_characterGenerator8x16[3332] = 8'h36;
assign _c_characterGenerator8x16[3333] = 8'h36;
assign _c_characterGenerator8x16[3334] = 8'h36;
assign _c_characterGenerator8x16[3335] = 8'hff;
assign _c_characterGenerator8x16[3336] = 8'h00;
assign _c_characterGenerator8x16[3337] = 8'h00;
assign _c_characterGenerator8x16[3338] = 8'h00;
assign _c_characterGenerator8x16[3339] = 8'h00;
assign _c_characterGenerator8x16[3340] = 8'h00;
assign _c_characterGenerator8x16[3341] = 8'h00;
assign _c_characterGenerator8x16[3342] = 8'h00;
assign _c_characterGenerator8x16[3343] = 8'h00;
assign _c_characterGenerator8x16[3344] = 8'h00;
assign _c_characterGenerator8x16[3345] = 8'h00;
assign _c_characterGenerator8x16[3346] = 8'h00;
assign _c_characterGenerator8x16[3347] = 8'h00;
assign _c_characterGenerator8x16[3348] = 8'h00;
assign _c_characterGenerator8x16[3349] = 8'hff;
assign _c_characterGenerator8x16[3350] = 8'h00;
assign _c_characterGenerator8x16[3351] = 8'hff;
assign _c_characterGenerator8x16[3352] = 8'h18;
assign _c_characterGenerator8x16[3353] = 8'h18;
assign _c_characterGenerator8x16[3354] = 8'h18;
assign _c_characterGenerator8x16[3355] = 8'h18;
assign _c_characterGenerator8x16[3356] = 8'h18;
assign _c_characterGenerator8x16[3357] = 8'h18;
assign _c_characterGenerator8x16[3358] = 8'h18;
assign _c_characterGenerator8x16[3359] = 8'h18;
assign _c_characterGenerator8x16[3360] = 8'h00;
assign _c_characterGenerator8x16[3361] = 8'h00;
assign _c_characterGenerator8x16[3362] = 8'h00;
assign _c_characterGenerator8x16[3363] = 8'h00;
assign _c_characterGenerator8x16[3364] = 8'h00;
assign _c_characterGenerator8x16[3365] = 8'h00;
assign _c_characterGenerator8x16[3366] = 8'h00;
assign _c_characterGenerator8x16[3367] = 8'hff;
assign _c_characterGenerator8x16[3368] = 8'h36;
assign _c_characterGenerator8x16[3369] = 8'h36;
assign _c_characterGenerator8x16[3370] = 8'h36;
assign _c_characterGenerator8x16[3371] = 8'h36;
assign _c_characterGenerator8x16[3372] = 8'h36;
assign _c_characterGenerator8x16[3373] = 8'h36;
assign _c_characterGenerator8x16[3374] = 8'h36;
assign _c_characterGenerator8x16[3375] = 8'h36;
assign _c_characterGenerator8x16[3376] = 8'h36;
assign _c_characterGenerator8x16[3377] = 8'h36;
assign _c_characterGenerator8x16[3378] = 8'h36;
assign _c_characterGenerator8x16[3379] = 8'h36;
assign _c_characterGenerator8x16[3380] = 8'h36;
assign _c_characterGenerator8x16[3381] = 8'h36;
assign _c_characterGenerator8x16[3382] = 8'h36;
assign _c_characterGenerator8x16[3383] = 8'h3f;
assign _c_characterGenerator8x16[3384] = 8'h00;
assign _c_characterGenerator8x16[3385] = 8'h00;
assign _c_characterGenerator8x16[3386] = 8'h00;
assign _c_characterGenerator8x16[3387] = 8'h00;
assign _c_characterGenerator8x16[3388] = 8'h00;
assign _c_characterGenerator8x16[3389] = 8'h00;
assign _c_characterGenerator8x16[3390] = 8'h00;
assign _c_characterGenerator8x16[3391] = 8'h00;
assign _c_characterGenerator8x16[3392] = 8'h18;
assign _c_characterGenerator8x16[3393] = 8'h18;
assign _c_characterGenerator8x16[3394] = 8'h18;
assign _c_characterGenerator8x16[3395] = 8'h18;
assign _c_characterGenerator8x16[3396] = 8'h18;
assign _c_characterGenerator8x16[3397] = 8'h1f;
assign _c_characterGenerator8x16[3398] = 8'h18;
assign _c_characterGenerator8x16[3399] = 8'h1f;
assign _c_characterGenerator8x16[3400] = 8'h00;
assign _c_characterGenerator8x16[3401] = 8'h00;
assign _c_characterGenerator8x16[3402] = 8'h00;
assign _c_characterGenerator8x16[3403] = 8'h00;
assign _c_characterGenerator8x16[3404] = 8'h00;
assign _c_characterGenerator8x16[3405] = 8'h00;
assign _c_characterGenerator8x16[3406] = 8'h00;
assign _c_characterGenerator8x16[3407] = 8'h00;
assign _c_characterGenerator8x16[3408] = 8'h00;
assign _c_characterGenerator8x16[3409] = 8'h00;
assign _c_characterGenerator8x16[3410] = 8'h00;
assign _c_characterGenerator8x16[3411] = 8'h00;
assign _c_characterGenerator8x16[3412] = 8'h00;
assign _c_characterGenerator8x16[3413] = 8'h1f;
assign _c_characterGenerator8x16[3414] = 8'h18;
assign _c_characterGenerator8x16[3415] = 8'h1f;
assign _c_characterGenerator8x16[3416] = 8'h18;
assign _c_characterGenerator8x16[3417] = 8'h18;
assign _c_characterGenerator8x16[3418] = 8'h18;
assign _c_characterGenerator8x16[3419] = 8'h18;
assign _c_characterGenerator8x16[3420] = 8'h18;
assign _c_characterGenerator8x16[3421] = 8'h18;
assign _c_characterGenerator8x16[3422] = 8'h18;
assign _c_characterGenerator8x16[3423] = 8'h18;
assign _c_characterGenerator8x16[3424] = 8'h00;
assign _c_characterGenerator8x16[3425] = 8'h00;
assign _c_characterGenerator8x16[3426] = 8'h00;
assign _c_characterGenerator8x16[3427] = 8'h00;
assign _c_characterGenerator8x16[3428] = 8'h00;
assign _c_characterGenerator8x16[3429] = 8'h00;
assign _c_characterGenerator8x16[3430] = 8'h00;
assign _c_characterGenerator8x16[3431] = 8'h3f;
assign _c_characterGenerator8x16[3432] = 8'h36;
assign _c_characterGenerator8x16[3433] = 8'h36;
assign _c_characterGenerator8x16[3434] = 8'h36;
assign _c_characterGenerator8x16[3435] = 8'h36;
assign _c_characterGenerator8x16[3436] = 8'h36;
assign _c_characterGenerator8x16[3437] = 8'h36;
assign _c_characterGenerator8x16[3438] = 8'h36;
assign _c_characterGenerator8x16[3439] = 8'h36;
assign _c_characterGenerator8x16[3440] = 8'h36;
assign _c_characterGenerator8x16[3441] = 8'h36;
assign _c_characterGenerator8x16[3442] = 8'h36;
assign _c_characterGenerator8x16[3443] = 8'h36;
assign _c_characterGenerator8x16[3444] = 8'h36;
assign _c_characterGenerator8x16[3445] = 8'h36;
assign _c_characterGenerator8x16[3446] = 8'h36;
assign _c_characterGenerator8x16[3447] = 8'hff;
assign _c_characterGenerator8x16[3448] = 8'h36;
assign _c_characterGenerator8x16[3449] = 8'h36;
assign _c_characterGenerator8x16[3450] = 8'h36;
assign _c_characterGenerator8x16[3451] = 8'h36;
assign _c_characterGenerator8x16[3452] = 8'h36;
assign _c_characterGenerator8x16[3453] = 8'h36;
assign _c_characterGenerator8x16[3454] = 8'h36;
assign _c_characterGenerator8x16[3455] = 8'h36;
assign _c_characterGenerator8x16[3456] = 8'h18;
assign _c_characterGenerator8x16[3457] = 8'h18;
assign _c_characterGenerator8x16[3458] = 8'h18;
assign _c_characterGenerator8x16[3459] = 8'h18;
assign _c_characterGenerator8x16[3460] = 8'h18;
assign _c_characterGenerator8x16[3461] = 8'hff;
assign _c_characterGenerator8x16[3462] = 8'h18;
assign _c_characterGenerator8x16[3463] = 8'hff;
assign _c_characterGenerator8x16[3464] = 8'h18;
assign _c_characterGenerator8x16[3465] = 8'h18;
assign _c_characterGenerator8x16[3466] = 8'h18;
assign _c_characterGenerator8x16[3467] = 8'h18;
assign _c_characterGenerator8x16[3468] = 8'h18;
assign _c_characterGenerator8x16[3469] = 8'h18;
assign _c_characterGenerator8x16[3470] = 8'h18;
assign _c_characterGenerator8x16[3471] = 8'h18;
assign _c_characterGenerator8x16[3472] = 8'h18;
assign _c_characterGenerator8x16[3473] = 8'h18;
assign _c_characterGenerator8x16[3474] = 8'h18;
assign _c_characterGenerator8x16[3475] = 8'h18;
assign _c_characterGenerator8x16[3476] = 8'h18;
assign _c_characterGenerator8x16[3477] = 8'h18;
assign _c_characterGenerator8x16[3478] = 8'h18;
assign _c_characterGenerator8x16[3479] = 8'hf8;
assign _c_characterGenerator8x16[3480] = 8'h00;
assign _c_characterGenerator8x16[3481] = 8'h00;
assign _c_characterGenerator8x16[3482] = 8'h00;
assign _c_characterGenerator8x16[3483] = 8'h00;
assign _c_characterGenerator8x16[3484] = 8'h00;
assign _c_characterGenerator8x16[3485] = 8'h00;
assign _c_characterGenerator8x16[3486] = 8'h00;
assign _c_characterGenerator8x16[3487] = 8'h00;
assign _c_characterGenerator8x16[3488] = 8'h00;
assign _c_characterGenerator8x16[3489] = 8'h00;
assign _c_characterGenerator8x16[3490] = 8'h00;
assign _c_characterGenerator8x16[3491] = 8'h00;
assign _c_characterGenerator8x16[3492] = 8'h00;
assign _c_characterGenerator8x16[3493] = 8'h00;
assign _c_characterGenerator8x16[3494] = 8'h00;
assign _c_characterGenerator8x16[3495] = 8'h1f;
assign _c_characterGenerator8x16[3496] = 8'h18;
assign _c_characterGenerator8x16[3497] = 8'h18;
assign _c_characterGenerator8x16[3498] = 8'h18;
assign _c_characterGenerator8x16[3499] = 8'h18;
assign _c_characterGenerator8x16[3500] = 8'h18;
assign _c_characterGenerator8x16[3501] = 8'h18;
assign _c_characterGenerator8x16[3502] = 8'h18;
assign _c_characterGenerator8x16[3503] = 8'h18;
assign _c_characterGenerator8x16[3504] = 8'hff;
assign _c_characterGenerator8x16[3505] = 8'hff;
assign _c_characterGenerator8x16[3506] = 8'hff;
assign _c_characterGenerator8x16[3507] = 8'hff;
assign _c_characterGenerator8x16[3508] = 8'hff;
assign _c_characterGenerator8x16[3509] = 8'hff;
assign _c_characterGenerator8x16[3510] = 8'hff;
assign _c_characterGenerator8x16[3511] = 8'hff;
assign _c_characterGenerator8x16[3512] = 8'hff;
assign _c_characterGenerator8x16[3513] = 8'hff;
assign _c_characterGenerator8x16[3514] = 8'hff;
assign _c_characterGenerator8x16[3515] = 8'hff;
assign _c_characterGenerator8x16[3516] = 8'hff;
assign _c_characterGenerator8x16[3517] = 8'hff;
assign _c_characterGenerator8x16[3518] = 8'hff;
assign _c_characterGenerator8x16[3519] = 8'hff;
assign _c_characterGenerator8x16[3520] = 8'h00;
assign _c_characterGenerator8x16[3521] = 8'h00;
assign _c_characterGenerator8x16[3522] = 8'h00;
assign _c_characterGenerator8x16[3523] = 8'h00;
assign _c_characterGenerator8x16[3524] = 8'h00;
assign _c_characterGenerator8x16[3525] = 8'h00;
assign _c_characterGenerator8x16[3526] = 8'h00;
assign _c_characterGenerator8x16[3527] = 8'hff;
assign _c_characterGenerator8x16[3528] = 8'hff;
assign _c_characterGenerator8x16[3529] = 8'hff;
assign _c_characterGenerator8x16[3530] = 8'hff;
assign _c_characterGenerator8x16[3531] = 8'hff;
assign _c_characterGenerator8x16[3532] = 8'hff;
assign _c_characterGenerator8x16[3533] = 8'hff;
assign _c_characterGenerator8x16[3534] = 8'hff;
assign _c_characterGenerator8x16[3535] = 8'hff;
assign _c_characterGenerator8x16[3536] = 8'hf0;
assign _c_characterGenerator8x16[3537] = 8'hf0;
assign _c_characterGenerator8x16[3538] = 8'hf0;
assign _c_characterGenerator8x16[3539] = 8'hf0;
assign _c_characterGenerator8x16[3540] = 8'hf0;
assign _c_characterGenerator8x16[3541] = 8'hf0;
assign _c_characterGenerator8x16[3542] = 8'hf0;
assign _c_characterGenerator8x16[3543] = 8'hf0;
assign _c_characterGenerator8x16[3544] = 8'hf0;
assign _c_characterGenerator8x16[3545] = 8'hf0;
assign _c_characterGenerator8x16[3546] = 8'hf0;
assign _c_characterGenerator8x16[3547] = 8'hf0;
assign _c_characterGenerator8x16[3548] = 8'hf0;
assign _c_characterGenerator8x16[3549] = 8'hf0;
assign _c_characterGenerator8x16[3550] = 8'hf0;
assign _c_characterGenerator8x16[3551] = 8'hf0;
assign _c_characterGenerator8x16[3552] = 8'h0f;
assign _c_characterGenerator8x16[3553] = 8'h0f;
assign _c_characterGenerator8x16[3554] = 8'h0f;
assign _c_characterGenerator8x16[3555] = 8'h0f;
assign _c_characterGenerator8x16[3556] = 8'h0f;
assign _c_characterGenerator8x16[3557] = 8'h0f;
assign _c_characterGenerator8x16[3558] = 8'h0f;
assign _c_characterGenerator8x16[3559] = 8'h0f;
assign _c_characterGenerator8x16[3560] = 8'h0f;
assign _c_characterGenerator8x16[3561] = 8'h0f;
assign _c_characterGenerator8x16[3562] = 8'h0f;
assign _c_characterGenerator8x16[3563] = 8'h0f;
assign _c_characterGenerator8x16[3564] = 8'h0f;
assign _c_characterGenerator8x16[3565] = 8'h0f;
assign _c_characterGenerator8x16[3566] = 8'h0f;
assign _c_characterGenerator8x16[3567] = 8'h0f;
assign _c_characterGenerator8x16[3568] = 8'hff;
assign _c_characterGenerator8x16[3569] = 8'hff;
assign _c_characterGenerator8x16[3570] = 8'hff;
assign _c_characterGenerator8x16[3571] = 8'hff;
assign _c_characterGenerator8x16[3572] = 8'hff;
assign _c_characterGenerator8x16[3573] = 8'hff;
assign _c_characterGenerator8x16[3574] = 8'hff;
assign _c_characterGenerator8x16[3575] = 8'h00;
assign _c_characterGenerator8x16[3576] = 8'h00;
assign _c_characterGenerator8x16[3577] = 8'h00;
assign _c_characterGenerator8x16[3578] = 8'h00;
assign _c_characterGenerator8x16[3579] = 8'h00;
assign _c_characterGenerator8x16[3580] = 8'h00;
assign _c_characterGenerator8x16[3581] = 8'h00;
assign _c_characterGenerator8x16[3582] = 8'h00;
assign _c_characterGenerator8x16[3583] = 8'h00;
assign _c_characterGenerator8x16[3584] = 8'h00;
assign _c_characterGenerator8x16[3585] = 8'h00;
assign _c_characterGenerator8x16[3586] = 8'h00;
assign _c_characterGenerator8x16[3587] = 8'h00;
assign _c_characterGenerator8x16[3588] = 8'h00;
assign _c_characterGenerator8x16[3589] = 8'h76;
assign _c_characterGenerator8x16[3590] = 8'hdc;
assign _c_characterGenerator8x16[3591] = 8'hd8;
assign _c_characterGenerator8x16[3592] = 8'hd8;
assign _c_characterGenerator8x16[3593] = 8'hd8;
assign _c_characterGenerator8x16[3594] = 8'hdc;
assign _c_characterGenerator8x16[3595] = 8'h76;
assign _c_characterGenerator8x16[3596] = 8'h00;
assign _c_characterGenerator8x16[3597] = 8'h00;
assign _c_characterGenerator8x16[3598] = 8'h00;
assign _c_characterGenerator8x16[3599] = 8'h00;
assign _c_characterGenerator8x16[3600] = 8'h00;
assign _c_characterGenerator8x16[3601] = 8'h00;
assign _c_characterGenerator8x16[3602] = 8'h78;
assign _c_characterGenerator8x16[3603] = 8'hcc;
assign _c_characterGenerator8x16[3604] = 8'hcc;
assign _c_characterGenerator8x16[3605] = 8'hcc;
assign _c_characterGenerator8x16[3606] = 8'hd8;
assign _c_characterGenerator8x16[3607] = 8'hcc;
assign _c_characterGenerator8x16[3608] = 8'hc6;
assign _c_characterGenerator8x16[3609] = 8'hc6;
assign _c_characterGenerator8x16[3610] = 8'hc6;
assign _c_characterGenerator8x16[3611] = 8'hcc;
assign _c_characterGenerator8x16[3612] = 8'h00;
assign _c_characterGenerator8x16[3613] = 8'h00;
assign _c_characterGenerator8x16[3614] = 8'h00;
assign _c_characterGenerator8x16[3615] = 8'h00;
assign _c_characterGenerator8x16[3616] = 8'h00;
assign _c_characterGenerator8x16[3617] = 8'h00;
assign _c_characterGenerator8x16[3618] = 8'hfe;
assign _c_characterGenerator8x16[3619] = 8'hc6;
assign _c_characterGenerator8x16[3620] = 8'hc6;
assign _c_characterGenerator8x16[3621] = 8'hc0;
assign _c_characterGenerator8x16[3622] = 8'hc0;
assign _c_characterGenerator8x16[3623] = 8'hc0;
assign _c_characterGenerator8x16[3624] = 8'hc0;
assign _c_characterGenerator8x16[3625] = 8'hc0;
assign _c_characterGenerator8x16[3626] = 8'hc0;
assign _c_characterGenerator8x16[3627] = 8'hc0;
assign _c_characterGenerator8x16[3628] = 8'h00;
assign _c_characterGenerator8x16[3629] = 8'h00;
assign _c_characterGenerator8x16[3630] = 8'h00;
assign _c_characterGenerator8x16[3631] = 8'h00;
assign _c_characterGenerator8x16[3632] = 8'h00;
assign _c_characterGenerator8x16[3633] = 8'h00;
assign _c_characterGenerator8x16[3634] = 8'h00;
assign _c_characterGenerator8x16[3635] = 8'h00;
assign _c_characterGenerator8x16[3636] = 8'hfe;
assign _c_characterGenerator8x16[3637] = 8'h6c;
assign _c_characterGenerator8x16[3638] = 8'h6c;
assign _c_characterGenerator8x16[3639] = 8'h6c;
assign _c_characterGenerator8x16[3640] = 8'h6c;
assign _c_characterGenerator8x16[3641] = 8'h6c;
assign _c_characterGenerator8x16[3642] = 8'h6c;
assign _c_characterGenerator8x16[3643] = 8'h6c;
assign _c_characterGenerator8x16[3644] = 8'h00;
assign _c_characterGenerator8x16[3645] = 8'h00;
assign _c_characterGenerator8x16[3646] = 8'h00;
assign _c_characterGenerator8x16[3647] = 8'h00;
assign _c_characterGenerator8x16[3648] = 8'h00;
assign _c_characterGenerator8x16[3649] = 8'h00;
assign _c_characterGenerator8x16[3650] = 8'h00;
assign _c_characterGenerator8x16[3651] = 8'hfe;
assign _c_characterGenerator8x16[3652] = 8'hc6;
assign _c_characterGenerator8x16[3653] = 8'h60;
assign _c_characterGenerator8x16[3654] = 8'h30;
assign _c_characterGenerator8x16[3655] = 8'h18;
assign _c_characterGenerator8x16[3656] = 8'h30;
assign _c_characterGenerator8x16[3657] = 8'h60;
assign _c_characterGenerator8x16[3658] = 8'hc6;
assign _c_characterGenerator8x16[3659] = 8'hfe;
assign _c_characterGenerator8x16[3660] = 8'h00;
assign _c_characterGenerator8x16[3661] = 8'h00;
assign _c_characterGenerator8x16[3662] = 8'h00;
assign _c_characterGenerator8x16[3663] = 8'h00;
assign _c_characterGenerator8x16[3664] = 8'h00;
assign _c_characterGenerator8x16[3665] = 8'h00;
assign _c_characterGenerator8x16[3666] = 8'h00;
assign _c_characterGenerator8x16[3667] = 8'h00;
assign _c_characterGenerator8x16[3668] = 8'h00;
assign _c_characterGenerator8x16[3669] = 8'h7e;
assign _c_characterGenerator8x16[3670] = 8'hd8;
assign _c_characterGenerator8x16[3671] = 8'hd8;
assign _c_characterGenerator8x16[3672] = 8'hd8;
assign _c_characterGenerator8x16[3673] = 8'hd8;
assign _c_characterGenerator8x16[3674] = 8'hd8;
assign _c_characterGenerator8x16[3675] = 8'h70;
assign _c_characterGenerator8x16[3676] = 8'h00;
assign _c_characterGenerator8x16[3677] = 8'h00;
assign _c_characterGenerator8x16[3678] = 8'h00;
assign _c_characterGenerator8x16[3679] = 8'h00;
assign _c_characterGenerator8x16[3680] = 8'h00;
assign _c_characterGenerator8x16[3681] = 8'h00;
assign _c_characterGenerator8x16[3682] = 8'h00;
assign _c_characterGenerator8x16[3683] = 8'h00;
assign _c_characterGenerator8x16[3684] = 8'h66;
assign _c_characterGenerator8x16[3685] = 8'h66;
assign _c_characterGenerator8x16[3686] = 8'h66;
assign _c_characterGenerator8x16[3687] = 8'h66;
assign _c_characterGenerator8x16[3688] = 8'h66;
assign _c_characterGenerator8x16[3689] = 8'h7c;
assign _c_characterGenerator8x16[3690] = 8'h60;
assign _c_characterGenerator8x16[3691] = 8'h60;
assign _c_characterGenerator8x16[3692] = 8'hc0;
assign _c_characterGenerator8x16[3693] = 8'h00;
assign _c_characterGenerator8x16[3694] = 8'h00;
assign _c_characterGenerator8x16[3695] = 8'h00;
assign _c_characterGenerator8x16[3696] = 8'h00;
assign _c_characterGenerator8x16[3697] = 8'h00;
assign _c_characterGenerator8x16[3698] = 8'h00;
assign _c_characterGenerator8x16[3699] = 8'h00;
assign _c_characterGenerator8x16[3700] = 8'h76;
assign _c_characterGenerator8x16[3701] = 8'hdc;
assign _c_characterGenerator8x16[3702] = 8'h18;
assign _c_characterGenerator8x16[3703] = 8'h18;
assign _c_characterGenerator8x16[3704] = 8'h18;
assign _c_characterGenerator8x16[3705] = 8'h18;
assign _c_characterGenerator8x16[3706] = 8'h18;
assign _c_characterGenerator8x16[3707] = 8'h18;
assign _c_characterGenerator8x16[3708] = 8'h00;
assign _c_characterGenerator8x16[3709] = 8'h00;
assign _c_characterGenerator8x16[3710] = 8'h00;
assign _c_characterGenerator8x16[3711] = 8'h00;
assign _c_characterGenerator8x16[3712] = 8'h00;
assign _c_characterGenerator8x16[3713] = 8'h00;
assign _c_characterGenerator8x16[3714] = 8'h00;
assign _c_characterGenerator8x16[3715] = 8'h7e;
assign _c_characterGenerator8x16[3716] = 8'h18;
assign _c_characterGenerator8x16[3717] = 8'h3c;
assign _c_characterGenerator8x16[3718] = 8'h66;
assign _c_characterGenerator8x16[3719] = 8'h66;
assign _c_characterGenerator8x16[3720] = 8'h66;
assign _c_characterGenerator8x16[3721] = 8'h3c;
assign _c_characterGenerator8x16[3722] = 8'h18;
assign _c_characterGenerator8x16[3723] = 8'h7e;
assign _c_characterGenerator8x16[3724] = 8'h00;
assign _c_characterGenerator8x16[3725] = 8'h00;
assign _c_characterGenerator8x16[3726] = 8'h00;
assign _c_characterGenerator8x16[3727] = 8'h00;
assign _c_characterGenerator8x16[3728] = 8'h00;
assign _c_characterGenerator8x16[3729] = 8'h00;
assign _c_characterGenerator8x16[3730] = 8'h00;
assign _c_characterGenerator8x16[3731] = 8'h38;
assign _c_characterGenerator8x16[3732] = 8'h6c;
assign _c_characterGenerator8x16[3733] = 8'hc6;
assign _c_characterGenerator8x16[3734] = 8'hc6;
assign _c_characterGenerator8x16[3735] = 8'hfe;
assign _c_characterGenerator8x16[3736] = 8'hc6;
assign _c_characterGenerator8x16[3737] = 8'hc6;
assign _c_characterGenerator8x16[3738] = 8'h6c;
assign _c_characterGenerator8x16[3739] = 8'h38;
assign _c_characterGenerator8x16[3740] = 8'h00;
assign _c_characterGenerator8x16[3741] = 8'h00;
assign _c_characterGenerator8x16[3742] = 8'h00;
assign _c_characterGenerator8x16[3743] = 8'h00;
assign _c_characterGenerator8x16[3744] = 8'h00;
assign _c_characterGenerator8x16[3745] = 8'h00;
assign _c_characterGenerator8x16[3746] = 8'h38;
assign _c_characterGenerator8x16[3747] = 8'h6c;
assign _c_characterGenerator8x16[3748] = 8'hc6;
assign _c_characterGenerator8x16[3749] = 8'hc6;
assign _c_characterGenerator8x16[3750] = 8'hc6;
assign _c_characterGenerator8x16[3751] = 8'h6c;
assign _c_characterGenerator8x16[3752] = 8'h6c;
assign _c_characterGenerator8x16[3753] = 8'h6c;
assign _c_characterGenerator8x16[3754] = 8'h6c;
assign _c_characterGenerator8x16[3755] = 8'hee;
assign _c_characterGenerator8x16[3756] = 8'h00;
assign _c_characterGenerator8x16[3757] = 8'h00;
assign _c_characterGenerator8x16[3758] = 8'h00;
assign _c_characterGenerator8x16[3759] = 8'h00;
assign _c_characterGenerator8x16[3760] = 8'h00;
assign _c_characterGenerator8x16[3761] = 8'h00;
assign _c_characterGenerator8x16[3762] = 8'h1e;
assign _c_characterGenerator8x16[3763] = 8'h30;
assign _c_characterGenerator8x16[3764] = 8'h18;
assign _c_characterGenerator8x16[3765] = 8'h0c;
assign _c_characterGenerator8x16[3766] = 8'h3e;
assign _c_characterGenerator8x16[3767] = 8'h66;
assign _c_characterGenerator8x16[3768] = 8'h66;
assign _c_characterGenerator8x16[3769] = 8'h66;
assign _c_characterGenerator8x16[3770] = 8'h66;
assign _c_characterGenerator8x16[3771] = 8'h3c;
assign _c_characterGenerator8x16[3772] = 8'h00;
assign _c_characterGenerator8x16[3773] = 8'h00;
assign _c_characterGenerator8x16[3774] = 8'h00;
assign _c_characterGenerator8x16[3775] = 8'h00;
assign _c_characterGenerator8x16[3776] = 8'h00;
assign _c_characterGenerator8x16[3777] = 8'h00;
assign _c_characterGenerator8x16[3778] = 8'h00;
assign _c_characterGenerator8x16[3779] = 8'h00;
assign _c_characterGenerator8x16[3780] = 8'h00;
assign _c_characterGenerator8x16[3781] = 8'h7e;
assign _c_characterGenerator8x16[3782] = 8'hdb;
assign _c_characterGenerator8x16[3783] = 8'hdb;
assign _c_characterGenerator8x16[3784] = 8'hdb;
assign _c_characterGenerator8x16[3785] = 8'h7e;
assign _c_characterGenerator8x16[3786] = 8'h00;
assign _c_characterGenerator8x16[3787] = 8'h00;
assign _c_characterGenerator8x16[3788] = 8'h00;
assign _c_characterGenerator8x16[3789] = 8'h00;
assign _c_characterGenerator8x16[3790] = 8'h00;
assign _c_characterGenerator8x16[3791] = 8'h00;
assign _c_characterGenerator8x16[3792] = 8'h00;
assign _c_characterGenerator8x16[3793] = 8'h00;
assign _c_characterGenerator8x16[3794] = 8'h00;
assign _c_characterGenerator8x16[3795] = 8'h03;
assign _c_characterGenerator8x16[3796] = 8'h06;
assign _c_characterGenerator8x16[3797] = 8'h7e;
assign _c_characterGenerator8x16[3798] = 8'hdb;
assign _c_characterGenerator8x16[3799] = 8'hdb;
assign _c_characterGenerator8x16[3800] = 8'hf3;
assign _c_characterGenerator8x16[3801] = 8'h7e;
assign _c_characterGenerator8x16[3802] = 8'h60;
assign _c_characterGenerator8x16[3803] = 8'hc0;
assign _c_characterGenerator8x16[3804] = 8'h00;
assign _c_characterGenerator8x16[3805] = 8'h00;
assign _c_characterGenerator8x16[3806] = 8'h00;
assign _c_characterGenerator8x16[3807] = 8'h00;
assign _c_characterGenerator8x16[3808] = 8'h00;
assign _c_characterGenerator8x16[3809] = 8'h00;
assign _c_characterGenerator8x16[3810] = 8'h1c;
assign _c_characterGenerator8x16[3811] = 8'h30;
assign _c_characterGenerator8x16[3812] = 8'h60;
assign _c_characterGenerator8x16[3813] = 8'h60;
assign _c_characterGenerator8x16[3814] = 8'h7c;
assign _c_characterGenerator8x16[3815] = 8'h60;
assign _c_characterGenerator8x16[3816] = 8'h60;
assign _c_characterGenerator8x16[3817] = 8'h60;
assign _c_characterGenerator8x16[3818] = 8'h30;
assign _c_characterGenerator8x16[3819] = 8'h1c;
assign _c_characterGenerator8x16[3820] = 8'h00;
assign _c_characterGenerator8x16[3821] = 8'h00;
assign _c_characterGenerator8x16[3822] = 8'h00;
assign _c_characterGenerator8x16[3823] = 8'h00;
assign _c_characterGenerator8x16[3824] = 8'h00;
assign _c_characterGenerator8x16[3825] = 8'h00;
assign _c_characterGenerator8x16[3826] = 8'h00;
assign _c_characterGenerator8x16[3827] = 8'h7c;
assign _c_characterGenerator8x16[3828] = 8'hc6;
assign _c_characterGenerator8x16[3829] = 8'hc6;
assign _c_characterGenerator8x16[3830] = 8'hc6;
assign _c_characterGenerator8x16[3831] = 8'hc6;
assign _c_characterGenerator8x16[3832] = 8'hc6;
assign _c_characterGenerator8x16[3833] = 8'hc6;
assign _c_characterGenerator8x16[3834] = 8'hc6;
assign _c_characterGenerator8x16[3835] = 8'hc6;
assign _c_characterGenerator8x16[3836] = 8'h00;
assign _c_characterGenerator8x16[3837] = 8'h00;
assign _c_characterGenerator8x16[3838] = 8'h00;
assign _c_characterGenerator8x16[3839] = 8'h00;
assign _c_characterGenerator8x16[3840] = 8'h00;
assign _c_characterGenerator8x16[3841] = 8'h00;
assign _c_characterGenerator8x16[3842] = 8'h00;
assign _c_characterGenerator8x16[3843] = 8'h00;
assign _c_characterGenerator8x16[3844] = 8'hfe;
assign _c_characterGenerator8x16[3845] = 8'h00;
assign _c_characterGenerator8x16[3846] = 8'h00;
assign _c_characterGenerator8x16[3847] = 8'hfe;
assign _c_characterGenerator8x16[3848] = 8'h00;
assign _c_characterGenerator8x16[3849] = 8'h00;
assign _c_characterGenerator8x16[3850] = 8'hfe;
assign _c_characterGenerator8x16[3851] = 8'h00;
assign _c_characterGenerator8x16[3852] = 8'h00;
assign _c_characterGenerator8x16[3853] = 8'h00;
assign _c_characterGenerator8x16[3854] = 8'h00;
assign _c_characterGenerator8x16[3855] = 8'h00;
assign _c_characterGenerator8x16[3856] = 8'h00;
assign _c_characterGenerator8x16[3857] = 8'h00;
assign _c_characterGenerator8x16[3858] = 8'h00;
assign _c_characterGenerator8x16[3859] = 8'h00;
assign _c_characterGenerator8x16[3860] = 8'h18;
assign _c_characterGenerator8x16[3861] = 8'h18;
assign _c_characterGenerator8x16[3862] = 8'h7e;
assign _c_characterGenerator8x16[3863] = 8'h18;
assign _c_characterGenerator8x16[3864] = 8'h18;
assign _c_characterGenerator8x16[3865] = 8'h00;
assign _c_characterGenerator8x16[3866] = 8'h00;
assign _c_characterGenerator8x16[3867] = 8'hff;
assign _c_characterGenerator8x16[3868] = 8'h00;
assign _c_characterGenerator8x16[3869] = 8'h00;
assign _c_characterGenerator8x16[3870] = 8'h00;
assign _c_characterGenerator8x16[3871] = 8'h00;
assign _c_characterGenerator8x16[3872] = 8'h00;
assign _c_characterGenerator8x16[3873] = 8'h00;
assign _c_characterGenerator8x16[3874] = 8'h00;
assign _c_characterGenerator8x16[3875] = 8'h30;
assign _c_characterGenerator8x16[3876] = 8'h18;
assign _c_characterGenerator8x16[3877] = 8'h0c;
assign _c_characterGenerator8x16[3878] = 8'h06;
assign _c_characterGenerator8x16[3879] = 8'h0c;
assign _c_characterGenerator8x16[3880] = 8'h18;
assign _c_characterGenerator8x16[3881] = 8'h30;
assign _c_characterGenerator8x16[3882] = 8'h00;
assign _c_characterGenerator8x16[3883] = 8'h7e;
assign _c_characterGenerator8x16[3884] = 8'h00;
assign _c_characterGenerator8x16[3885] = 8'h00;
assign _c_characterGenerator8x16[3886] = 8'h00;
assign _c_characterGenerator8x16[3887] = 8'h00;
assign _c_characterGenerator8x16[3888] = 8'h00;
assign _c_characterGenerator8x16[3889] = 8'h00;
assign _c_characterGenerator8x16[3890] = 8'h00;
assign _c_characterGenerator8x16[3891] = 8'h0c;
assign _c_characterGenerator8x16[3892] = 8'h18;
assign _c_characterGenerator8x16[3893] = 8'h30;
assign _c_characterGenerator8x16[3894] = 8'h60;
assign _c_characterGenerator8x16[3895] = 8'h30;
assign _c_characterGenerator8x16[3896] = 8'h18;
assign _c_characterGenerator8x16[3897] = 8'h0c;
assign _c_characterGenerator8x16[3898] = 8'h00;
assign _c_characterGenerator8x16[3899] = 8'h7e;
assign _c_characterGenerator8x16[3900] = 8'h00;
assign _c_characterGenerator8x16[3901] = 8'h00;
assign _c_characterGenerator8x16[3902] = 8'h00;
assign _c_characterGenerator8x16[3903] = 8'h00;
assign _c_characterGenerator8x16[3904] = 8'h00;
assign _c_characterGenerator8x16[3905] = 8'h00;
assign _c_characterGenerator8x16[3906] = 8'h0e;
assign _c_characterGenerator8x16[3907] = 8'h1b;
assign _c_characterGenerator8x16[3908] = 8'h1b;
assign _c_characterGenerator8x16[3909] = 8'h18;
assign _c_characterGenerator8x16[3910] = 8'h18;
assign _c_characterGenerator8x16[3911] = 8'h18;
assign _c_characterGenerator8x16[3912] = 8'h18;
assign _c_characterGenerator8x16[3913] = 8'h18;
assign _c_characterGenerator8x16[3914] = 8'h18;
assign _c_characterGenerator8x16[3915] = 8'h18;
assign _c_characterGenerator8x16[3916] = 8'h18;
assign _c_characterGenerator8x16[3917] = 8'h18;
assign _c_characterGenerator8x16[3918] = 8'h18;
assign _c_characterGenerator8x16[3919] = 8'h18;
assign _c_characterGenerator8x16[3920] = 8'h18;
assign _c_characterGenerator8x16[3921] = 8'h18;
assign _c_characterGenerator8x16[3922] = 8'h18;
assign _c_characterGenerator8x16[3923] = 8'h18;
assign _c_characterGenerator8x16[3924] = 8'h18;
assign _c_characterGenerator8x16[3925] = 8'h18;
assign _c_characterGenerator8x16[3926] = 8'h18;
assign _c_characterGenerator8x16[3927] = 8'h18;
assign _c_characterGenerator8x16[3928] = 8'hd8;
assign _c_characterGenerator8x16[3929] = 8'hd8;
assign _c_characterGenerator8x16[3930] = 8'hd8;
assign _c_characterGenerator8x16[3931] = 8'h70;
assign _c_characterGenerator8x16[3932] = 8'h00;
assign _c_characterGenerator8x16[3933] = 8'h00;
assign _c_characterGenerator8x16[3934] = 8'h00;
assign _c_characterGenerator8x16[3935] = 8'h00;
assign _c_characterGenerator8x16[3936] = 8'h00;
assign _c_characterGenerator8x16[3937] = 8'h00;
assign _c_characterGenerator8x16[3938] = 8'h00;
assign _c_characterGenerator8x16[3939] = 8'h00;
assign _c_characterGenerator8x16[3940] = 8'h18;
assign _c_characterGenerator8x16[3941] = 8'h18;
assign _c_characterGenerator8x16[3942] = 8'h00;
assign _c_characterGenerator8x16[3943] = 8'h7e;
assign _c_characterGenerator8x16[3944] = 8'h00;
assign _c_characterGenerator8x16[3945] = 8'h18;
assign _c_characterGenerator8x16[3946] = 8'h18;
assign _c_characterGenerator8x16[3947] = 8'h00;
assign _c_characterGenerator8x16[3948] = 8'h00;
assign _c_characterGenerator8x16[3949] = 8'h00;
assign _c_characterGenerator8x16[3950] = 8'h00;
assign _c_characterGenerator8x16[3951] = 8'h00;
assign _c_characterGenerator8x16[3952] = 8'h00;
assign _c_characterGenerator8x16[3953] = 8'h00;
assign _c_characterGenerator8x16[3954] = 8'h00;
assign _c_characterGenerator8x16[3955] = 8'h00;
assign _c_characterGenerator8x16[3956] = 8'h00;
assign _c_characterGenerator8x16[3957] = 8'h76;
assign _c_characterGenerator8x16[3958] = 8'hdc;
assign _c_characterGenerator8x16[3959] = 8'h00;
assign _c_characterGenerator8x16[3960] = 8'h76;
assign _c_characterGenerator8x16[3961] = 8'hdc;
assign _c_characterGenerator8x16[3962] = 8'h00;
assign _c_characterGenerator8x16[3963] = 8'h00;
assign _c_characterGenerator8x16[3964] = 8'h00;
assign _c_characterGenerator8x16[3965] = 8'h00;
assign _c_characterGenerator8x16[3966] = 8'h00;
assign _c_characterGenerator8x16[3967] = 8'h00;
assign _c_characterGenerator8x16[3968] = 8'h00;
assign _c_characterGenerator8x16[3969] = 8'h38;
assign _c_characterGenerator8x16[3970] = 8'h6c;
assign _c_characterGenerator8x16[3971] = 8'h6c;
assign _c_characterGenerator8x16[3972] = 8'h38;
assign _c_characterGenerator8x16[3973] = 8'h00;
assign _c_characterGenerator8x16[3974] = 8'h00;
assign _c_characterGenerator8x16[3975] = 8'h00;
assign _c_characterGenerator8x16[3976] = 8'h00;
assign _c_characterGenerator8x16[3977] = 8'h00;
assign _c_characterGenerator8x16[3978] = 8'h00;
assign _c_characterGenerator8x16[3979] = 8'h00;
assign _c_characterGenerator8x16[3980] = 8'h00;
assign _c_characterGenerator8x16[3981] = 8'h00;
assign _c_characterGenerator8x16[3982] = 8'h00;
assign _c_characterGenerator8x16[3983] = 8'h00;
assign _c_characterGenerator8x16[3984] = 8'h00;
assign _c_characterGenerator8x16[3985] = 8'h00;
assign _c_characterGenerator8x16[3986] = 8'h00;
assign _c_characterGenerator8x16[3987] = 8'h00;
assign _c_characterGenerator8x16[3988] = 8'h00;
assign _c_characterGenerator8x16[3989] = 8'h00;
assign _c_characterGenerator8x16[3990] = 8'h00;
assign _c_characterGenerator8x16[3991] = 8'h18;
assign _c_characterGenerator8x16[3992] = 8'h18;
assign _c_characterGenerator8x16[3993] = 8'h00;
assign _c_characterGenerator8x16[3994] = 8'h00;
assign _c_characterGenerator8x16[3995] = 8'h00;
assign _c_characterGenerator8x16[3996] = 8'h00;
assign _c_characterGenerator8x16[3997] = 8'h00;
assign _c_characterGenerator8x16[3998] = 8'h00;
assign _c_characterGenerator8x16[3999] = 8'h00;
assign _c_characterGenerator8x16[4000] = 8'h00;
assign _c_characterGenerator8x16[4001] = 8'h00;
assign _c_characterGenerator8x16[4002] = 8'h00;
assign _c_characterGenerator8x16[4003] = 8'h00;
assign _c_characterGenerator8x16[4004] = 8'h00;
assign _c_characterGenerator8x16[4005] = 8'h00;
assign _c_characterGenerator8x16[4006] = 8'h00;
assign _c_characterGenerator8x16[4007] = 8'h00;
assign _c_characterGenerator8x16[4008] = 8'h18;
assign _c_characterGenerator8x16[4009] = 8'h00;
assign _c_characterGenerator8x16[4010] = 8'h00;
assign _c_characterGenerator8x16[4011] = 8'h00;
assign _c_characterGenerator8x16[4012] = 8'h00;
assign _c_characterGenerator8x16[4013] = 8'h00;
assign _c_characterGenerator8x16[4014] = 8'h00;
assign _c_characterGenerator8x16[4015] = 8'h00;
assign _c_characterGenerator8x16[4016] = 8'h00;
assign _c_characterGenerator8x16[4017] = 8'h0f;
assign _c_characterGenerator8x16[4018] = 8'h0c;
assign _c_characterGenerator8x16[4019] = 8'h0c;
assign _c_characterGenerator8x16[4020] = 8'h0c;
assign _c_characterGenerator8x16[4021] = 8'h0c;
assign _c_characterGenerator8x16[4022] = 8'h0c;
assign _c_characterGenerator8x16[4023] = 8'hec;
assign _c_characterGenerator8x16[4024] = 8'h6c;
assign _c_characterGenerator8x16[4025] = 8'h6c;
assign _c_characterGenerator8x16[4026] = 8'h3c;
assign _c_characterGenerator8x16[4027] = 8'h1c;
assign _c_characterGenerator8x16[4028] = 8'h00;
assign _c_characterGenerator8x16[4029] = 8'h00;
assign _c_characterGenerator8x16[4030] = 8'h00;
assign _c_characterGenerator8x16[4031] = 8'h00;
assign _c_characterGenerator8x16[4032] = 8'h00;
assign _c_characterGenerator8x16[4033] = 8'hd8;
assign _c_characterGenerator8x16[4034] = 8'h6c;
assign _c_characterGenerator8x16[4035] = 8'h6c;
assign _c_characterGenerator8x16[4036] = 8'h6c;
assign _c_characterGenerator8x16[4037] = 8'h6c;
assign _c_characterGenerator8x16[4038] = 8'h6c;
assign _c_characterGenerator8x16[4039] = 8'h00;
assign _c_characterGenerator8x16[4040] = 8'h00;
assign _c_characterGenerator8x16[4041] = 8'h00;
assign _c_characterGenerator8x16[4042] = 8'h00;
assign _c_characterGenerator8x16[4043] = 8'h00;
assign _c_characterGenerator8x16[4044] = 8'h00;
assign _c_characterGenerator8x16[4045] = 8'h00;
assign _c_characterGenerator8x16[4046] = 8'h00;
assign _c_characterGenerator8x16[4047] = 8'h00;
assign _c_characterGenerator8x16[4048] = 8'h00;
assign _c_characterGenerator8x16[4049] = 8'h70;
assign _c_characterGenerator8x16[4050] = 8'hd8;
assign _c_characterGenerator8x16[4051] = 8'h30;
assign _c_characterGenerator8x16[4052] = 8'h60;
assign _c_characterGenerator8x16[4053] = 8'hc8;
assign _c_characterGenerator8x16[4054] = 8'hf8;
assign _c_characterGenerator8x16[4055] = 8'h00;
assign _c_characterGenerator8x16[4056] = 8'h00;
assign _c_characterGenerator8x16[4057] = 8'h00;
assign _c_characterGenerator8x16[4058] = 8'h00;
assign _c_characterGenerator8x16[4059] = 8'h00;
assign _c_characterGenerator8x16[4060] = 8'h00;
assign _c_characterGenerator8x16[4061] = 8'h00;
assign _c_characterGenerator8x16[4062] = 8'h00;
assign _c_characterGenerator8x16[4063] = 8'h00;
assign _c_characterGenerator8x16[4064] = 8'h00;
assign _c_characterGenerator8x16[4065] = 8'h00;
assign _c_characterGenerator8x16[4066] = 8'h00;
assign _c_characterGenerator8x16[4067] = 8'h00;
assign _c_characterGenerator8x16[4068] = 8'h7c;
assign _c_characterGenerator8x16[4069] = 8'h7c;
assign _c_characterGenerator8x16[4070] = 8'h7c;
assign _c_characterGenerator8x16[4071] = 8'h7c;
assign _c_characterGenerator8x16[4072] = 8'h7c;
assign _c_characterGenerator8x16[4073] = 8'h7c;
assign _c_characterGenerator8x16[4074] = 8'h7c;
assign _c_characterGenerator8x16[4075] = 8'h00;
assign _c_characterGenerator8x16[4076] = 8'h00;
assign _c_characterGenerator8x16[4077] = 8'h00;
assign _c_characterGenerator8x16[4078] = 8'h00;
assign _c_characterGenerator8x16[4079] = 8'h00;
assign _c_characterGenerator8x16[4080] = 8'h00;
assign _c_characterGenerator8x16[4081] = 8'h00;
assign _c_characterGenerator8x16[4082] = 8'h00;
assign _c_characterGenerator8x16[4083] = 8'h00;
assign _c_characterGenerator8x16[4084] = 8'h00;
assign _c_characterGenerator8x16[4085] = 8'h00;
assign _c_characterGenerator8x16[4086] = 8'h00;
assign _c_characterGenerator8x16[4087] = 8'h00;
assign _c_characterGenerator8x16[4088] = 8'h00;
assign _c_characterGenerator8x16[4089] = 8'h00;
assign _c_characterGenerator8x16[4090] = 8'h00;
assign _c_characterGenerator8x16[4091] = 8'h00;
assign _c_characterGenerator8x16[4092] = 8'h00;
assign _c_characterGenerator8x16[4093] = 8'h00;
assign _c_characterGenerator8x16[4094] = 8'h00;
assign _c_characterGenerator8x16[4095] = 8'h00;
wire  [7:0] _c_characterGenerator8x8[2047:0];
assign _c_characterGenerator8x8[0] = 8'h00;
assign _c_characterGenerator8x8[1] = 8'h00;
assign _c_characterGenerator8x8[2] = 8'h00;
assign _c_characterGenerator8x8[3] = 8'h00;
assign _c_characterGenerator8x8[4] = 8'h00;
assign _c_characterGenerator8x8[5] = 8'h00;
assign _c_characterGenerator8x8[6] = 8'h00;
assign _c_characterGenerator8x8[7] = 8'h00;
assign _c_characterGenerator8x8[8] = 8'h7e;
assign _c_characterGenerator8x8[9] = 8'h81;
assign _c_characterGenerator8x8[10] = 8'ha5;
assign _c_characterGenerator8x8[11] = 8'h81;
assign _c_characterGenerator8x8[12] = 8'hbd;
assign _c_characterGenerator8x8[13] = 8'h99;
assign _c_characterGenerator8x8[14] = 8'h81;
assign _c_characterGenerator8x8[15] = 8'h7e;
assign _c_characterGenerator8x8[16] = 8'h7e;
assign _c_characterGenerator8x8[17] = 8'hff;
assign _c_characterGenerator8x8[18] = 8'hdb;
assign _c_characterGenerator8x8[19] = 8'hff;
assign _c_characterGenerator8x8[20] = 8'hc3;
assign _c_characterGenerator8x8[21] = 8'he7;
assign _c_characterGenerator8x8[22] = 8'hff;
assign _c_characterGenerator8x8[23] = 8'h7e;
assign _c_characterGenerator8x8[24] = 8'h6c;
assign _c_characterGenerator8x8[25] = 8'hfe;
assign _c_characterGenerator8x8[26] = 8'hfe;
assign _c_characterGenerator8x8[27] = 8'hfe;
assign _c_characterGenerator8x8[28] = 8'h7c;
assign _c_characterGenerator8x8[29] = 8'h38;
assign _c_characterGenerator8x8[30] = 8'h10;
assign _c_characterGenerator8x8[31] = 8'h00;
assign _c_characterGenerator8x8[32] = 8'h10;
assign _c_characterGenerator8x8[33] = 8'h38;
assign _c_characterGenerator8x8[34] = 8'h7c;
assign _c_characterGenerator8x8[35] = 8'hfe;
assign _c_characterGenerator8x8[36] = 8'h7c;
assign _c_characterGenerator8x8[37] = 8'h38;
assign _c_characterGenerator8x8[38] = 8'h10;
assign _c_characterGenerator8x8[39] = 8'h00;
assign _c_characterGenerator8x8[40] = 8'h38;
assign _c_characterGenerator8x8[41] = 8'h7c;
assign _c_characterGenerator8x8[42] = 8'h38;
assign _c_characterGenerator8x8[43] = 8'hfe;
assign _c_characterGenerator8x8[44] = 8'hfe;
assign _c_characterGenerator8x8[45] = 8'h7c;
assign _c_characterGenerator8x8[46] = 8'h38;
assign _c_characterGenerator8x8[47] = 8'h7c;
assign _c_characterGenerator8x8[48] = 8'h10;
assign _c_characterGenerator8x8[49] = 8'h10;
assign _c_characterGenerator8x8[50] = 8'h38;
assign _c_characterGenerator8x8[51] = 8'h7c;
assign _c_characterGenerator8x8[52] = 8'hfe;
assign _c_characterGenerator8x8[53] = 8'h7c;
assign _c_characterGenerator8x8[54] = 8'h38;
assign _c_characterGenerator8x8[55] = 8'h7c;
assign _c_characterGenerator8x8[56] = 8'h00;
assign _c_characterGenerator8x8[57] = 8'h00;
assign _c_characterGenerator8x8[58] = 8'h18;
assign _c_characterGenerator8x8[59] = 8'h3c;
assign _c_characterGenerator8x8[60] = 8'h3c;
assign _c_characterGenerator8x8[61] = 8'h18;
assign _c_characterGenerator8x8[62] = 8'h00;
assign _c_characterGenerator8x8[63] = 8'h00;
assign _c_characterGenerator8x8[64] = 8'hff;
assign _c_characterGenerator8x8[65] = 8'hff;
assign _c_characterGenerator8x8[66] = 8'he7;
assign _c_characterGenerator8x8[67] = 8'hc3;
assign _c_characterGenerator8x8[68] = 8'hc3;
assign _c_characterGenerator8x8[69] = 8'he7;
assign _c_characterGenerator8x8[70] = 8'hff;
assign _c_characterGenerator8x8[71] = 8'hff;
assign _c_characterGenerator8x8[72] = 8'h00;
assign _c_characterGenerator8x8[73] = 8'h3c;
assign _c_characterGenerator8x8[74] = 8'h66;
assign _c_characterGenerator8x8[75] = 8'h42;
assign _c_characterGenerator8x8[76] = 8'h42;
assign _c_characterGenerator8x8[77] = 8'h66;
assign _c_characterGenerator8x8[78] = 8'h3c;
assign _c_characterGenerator8x8[79] = 8'h00;
assign _c_characterGenerator8x8[80] = 8'hff;
assign _c_characterGenerator8x8[81] = 8'hc3;
assign _c_characterGenerator8x8[82] = 8'h99;
assign _c_characterGenerator8x8[83] = 8'hbd;
assign _c_characterGenerator8x8[84] = 8'hbd;
assign _c_characterGenerator8x8[85] = 8'h99;
assign _c_characterGenerator8x8[86] = 8'hc3;
assign _c_characterGenerator8x8[87] = 8'hff;
assign _c_characterGenerator8x8[88] = 8'h0f;
assign _c_characterGenerator8x8[89] = 8'h07;
assign _c_characterGenerator8x8[90] = 8'h0f;
assign _c_characterGenerator8x8[91] = 8'h7d;
assign _c_characterGenerator8x8[92] = 8'hcc;
assign _c_characterGenerator8x8[93] = 8'hcc;
assign _c_characterGenerator8x8[94] = 8'hcc;
assign _c_characterGenerator8x8[95] = 8'h78;
assign _c_characterGenerator8x8[96] = 8'h3c;
assign _c_characterGenerator8x8[97] = 8'h66;
assign _c_characterGenerator8x8[98] = 8'h66;
assign _c_characterGenerator8x8[99] = 8'h66;
assign _c_characterGenerator8x8[100] = 8'h3c;
assign _c_characterGenerator8x8[101] = 8'h18;
assign _c_characterGenerator8x8[102] = 8'h7e;
assign _c_characterGenerator8x8[103] = 8'h18;
assign _c_characterGenerator8x8[104] = 8'h3f;
assign _c_characterGenerator8x8[105] = 8'h33;
assign _c_characterGenerator8x8[106] = 8'h3f;
assign _c_characterGenerator8x8[107] = 8'h30;
assign _c_characterGenerator8x8[108] = 8'h30;
assign _c_characterGenerator8x8[109] = 8'h70;
assign _c_characterGenerator8x8[110] = 8'hf0;
assign _c_characterGenerator8x8[111] = 8'he0;
assign _c_characterGenerator8x8[112] = 8'h7f;
assign _c_characterGenerator8x8[113] = 8'h63;
assign _c_characterGenerator8x8[114] = 8'h7f;
assign _c_characterGenerator8x8[115] = 8'h63;
assign _c_characterGenerator8x8[116] = 8'h63;
assign _c_characterGenerator8x8[117] = 8'h67;
assign _c_characterGenerator8x8[118] = 8'he6;
assign _c_characterGenerator8x8[119] = 8'hc0;
assign _c_characterGenerator8x8[120] = 8'h99;
assign _c_characterGenerator8x8[121] = 8'h5a;
assign _c_characterGenerator8x8[122] = 8'h3c;
assign _c_characterGenerator8x8[123] = 8'he7;
assign _c_characterGenerator8x8[124] = 8'he7;
assign _c_characterGenerator8x8[125] = 8'h3c;
assign _c_characterGenerator8x8[126] = 8'h5a;
assign _c_characterGenerator8x8[127] = 8'h99;
assign _c_characterGenerator8x8[128] = 8'h80;
assign _c_characterGenerator8x8[129] = 8'he0;
assign _c_characterGenerator8x8[130] = 8'hf8;
assign _c_characterGenerator8x8[131] = 8'hfe;
assign _c_characterGenerator8x8[132] = 8'hf8;
assign _c_characterGenerator8x8[133] = 8'he0;
assign _c_characterGenerator8x8[134] = 8'h80;
assign _c_characterGenerator8x8[135] = 8'h00;
assign _c_characterGenerator8x8[136] = 8'h02;
assign _c_characterGenerator8x8[137] = 8'h0e;
assign _c_characterGenerator8x8[138] = 8'h3e;
assign _c_characterGenerator8x8[139] = 8'hfe;
assign _c_characterGenerator8x8[140] = 8'h3e;
assign _c_characterGenerator8x8[141] = 8'h0e;
assign _c_characterGenerator8x8[142] = 8'h02;
assign _c_characterGenerator8x8[143] = 8'h00;
assign _c_characterGenerator8x8[144] = 8'h18;
assign _c_characterGenerator8x8[145] = 8'h3c;
assign _c_characterGenerator8x8[146] = 8'h7e;
assign _c_characterGenerator8x8[147] = 8'h18;
assign _c_characterGenerator8x8[148] = 8'h18;
assign _c_characterGenerator8x8[149] = 8'h7e;
assign _c_characterGenerator8x8[150] = 8'h3c;
assign _c_characterGenerator8x8[151] = 8'h18;
assign _c_characterGenerator8x8[152] = 8'h66;
assign _c_characterGenerator8x8[153] = 8'h66;
assign _c_characterGenerator8x8[154] = 8'h66;
assign _c_characterGenerator8x8[155] = 8'h66;
assign _c_characterGenerator8x8[156] = 8'h66;
assign _c_characterGenerator8x8[157] = 8'h00;
assign _c_characterGenerator8x8[158] = 8'h66;
assign _c_characterGenerator8x8[159] = 8'h00;
assign _c_characterGenerator8x8[160] = 8'h7f;
assign _c_characterGenerator8x8[161] = 8'hdb;
assign _c_characterGenerator8x8[162] = 8'hdb;
assign _c_characterGenerator8x8[163] = 8'h7b;
assign _c_characterGenerator8x8[164] = 8'h1b;
assign _c_characterGenerator8x8[165] = 8'h1b;
assign _c_characterGenerator8x8[166] = 8'h1b;
assign _c_characterGenerator8x8[167] = 8'h00;
assign _c_characterGenerator8x8[168] = 8'h3e;
assign _c_characterGenerator8x8[169] = 8'h63;
assign _c_characterGenerator8x8[170] = 8'h38;
assign _c_characterGenerator8x8[171] = 8'h6c;
assign _c_characterGenerator8x8[172] = 8'h6c;
assign _c_characterGenerator8x8[173] = 8'h38;
assign _c_characterGenerator8x8[174] = 8'hcc;
assign _c_characterGenerator8x8[175] = 8'h78;
assign _c_characterGenerator8x8[176] = 8'h00;
assign _c_characterGenerator8x8[177] = 8'h00;
assign _c_characterGenerator8x8[178] = 8'h00;
assign _c_characterGenerator8x8[179] = 8'h00;
assign _c_characterGenerator8x8[180] = 8'h7e;
assign _c_characterGenerator8x8[181] = 8'h7e;
assign _c_characterGenerator8x8[182] = 8'h7e;
assign _c_characterGenerator8x8[183] = 8'h00;
assign _c_characterGenerator8x8[184] = 8'h18;
assign _c_characterGenerator8x8[185] = 8'h3c;
assign _c_characterGenerator8x8[186] = 8'h7e;
assign _c_characterGenerator8x8[187] = 8'h18;
assign _c_characterGenerator8x8[188] = 8'h7e;
assign _c_characterGenerator8x8[189] = 8'h3c;
assign _c_characterGenerator8x8[190] = 8'h18;
assign _c_characterGenerator8x8[191] = 8'hff;
assign _c_characterGenerator8x8[192] = 8'h18;
assign _c_characterGenerator8x8[193] = 8'h3c;
assign _c_characterGenerator8x8[194] = 8'h7e;
assign _c_characterGenerator8x8[195] = 8'h18;
assign _c_characterGenerator8x8[196] = 8'h18;
assign _c_characterGenerator8x8[197] = 8'h18;
assign _c_characterGenerator8x8[198] = 8'h18;
assign _c_characterGenerator8x8[199] = 8'h00;
assign _c_characterGenerator8x8[200] = 8'h18;
assign _c_characterGenerator8x8[201] = 8'h18;
assign _c_characterGenerator8x8[202] = 8'h18;
assign _c_characterGenerator8x8[203] = 8'h18;
assign _c_characterGenerator8x8[204] = 8'h7e;
assign _c_characterGenerator8x8[205] = 8'h3c;
assign _c_characterGenerator8x8[206] = 8'h18;
assign _c_characterGenerator8x8[207] = 8'h00;
assign _c_characterGenerator8x8[208] = 8'h00;
assign _c_characterGenerator8x8[209] = 8'h18;
assign _c_characterGenerator8x8[210] = 8'h0c;
assign _c_characterGenerator8x8[211] = 8'hfe;
assign _c_characterGenerator8x8[212] = 8'h0c;
assign _c_characterGenerator8x8[213] = 8'h18;
assign _c_characterGenerator8x8[214] = 8'h00;
assign _c_characterGenerator8x8[215] = 8'h00;
assign _c_characterGenerator8x8[216] = 8'h00;
assign _c_characterGenerator8x8[217] = 8'h30;
assign _c_characterGenerator8x8[218] = 8'h60;
assign _c_characterGenerator8x8[219] = 8'hfe;
assign _c_characterGenerator8x8[220] = 8'h60;
assign _c_characterGenerator8x8[221] = 8'h30;
assign _c_characterGenerator8x8[222] = 8'h00;
assign _c_characterGenerator8x8[223] = 8'h00;
assign _c_characterGenerator8x8[224] = 8'h00;
assign _c_characterGenerator8x8[225] = 8'h00;
assign _c_characterGenerator8x8[226] = 8'hc0;
assign _c_characterGenerator8x8[227] = 8'hc0;
assign _c_characterGenerator8x8[228] = 8'hc0;
assign _c_characterGenerator8x8[229] = 8'hfe;
assign _c_characterGenerator8x8[230] = 8'h00;
assign _c_characterGenerator8x8[231] = 8'h00;
assign _c_characterGenerator8x8[232] = 8'h00;
assign _c_characterGenerator8x8[233] = 8'h24;
assign _c_characterGenerator8x8[234] = 8'h66;
assign _c_characterGenerator8x8[235] = 8'hff;
assign _c_characterGenerator8x8[236] = 8'h66;
assign _c_characterGenerator8x8[237] = 8'h24;
assign _c_characterGenerator8x8[238] = 8'h00;
assign _c_characterGenerator8x8[239] = 8'h00;
assign _c_characterGenerator8x8[240] = 8'h00;
assign _c_characterGenerator8x8[241] = 8'h18;
assign _c_characterGenerator8x8[242] = 8'h3c;
assign _c_characterGenerator8x8[243] = 8'h7e;
assign _c_characterGenerator8x8[244] = 8'hff;
assign _c_characterGenerator8x8[245] = 8'hff;
assign _c_characterGenerator8x8[246] = 8'h00;
assign _c_characterGenerator8x8[247] = 8'h00;
assign _c_characterGenerator8x8[248] = 8'h00;
assign _c_characterGenerator8x8[249] = 8'hff;
assign _c_characterGenerator8x8[250] = 8'hff;
assign _c_characterGenerator8x8[251] = 8'h7e;
assign _c_characterGenerator8x8[252] = 8'h3c;
assign _c_characterGenerator8x8[253] = 8'h18;
assign _c_characterGenerator8x8[254] = 8'h00;
assign _c_characterGenerator8x8[255] = 8'h00;
assign _c_characterGenerator8x8[256] = 8'h00;
assign _c_characterGenerator8x8[257] = 8'h00;
assign _c_characterGenerator8x8[258] = 8'h00;
assign _c_characterGenerator8x8[259] = 8'h00;
assign _c_characterGenerator8x8[260] = 8'h00;
assign _c_characterGenerator8x8[261] = 8'h00;
assign _c_characterGenerator8x8[262] = 8'h00;
assign _c_characterGenerator8x8[263] = 8'h00;
assign _c_characterGenerator8x8[264] = 8'h30;
assign _c_characterGenerator8x8[265] = 8'h78;
assign _c_characterGenerator8x8[266] = 8'h78;
assign _c_characterGenerator8x8[267] = 8'h30;
assign _c_characterGenerator8x8[268] = 8'h30;
assign _c_characterGenerator8x8[269] = 8'h00;
assign _c_characterGenerator8x8[270] = 8'h30;
assign _c_characterGenerator8x8[271] = 8'h00;
assign _c_characterGenerator8x8[272] = 8'h6c;
assign _c_characterGenerator8x8[273] = 8'h6c;
assign _c_characterGenerator8x8[274] = 8'h6c;
assign _c_characterGenerator8x8[275] = 8'h00;
assign _c_characterGenerator8x8[276] = 8'h00;
assign _c_characterGenerator8x8[277] = 8'h00;
assign _c_characterGenerator8x8[278] = 8'h00;
assign _c_characterGenerator8x8[279] = 8'h00;
assign _c_characterGenerator8x8[280] = 8'h6c;
assign _c_characterGenerator8x8[281] = 8'h6c;
assign _c_characterGenerator8x8[282] = 8'hfe;
assign _c_characterGenerator8x8[283] = 8'h6c;
assign _c_characterGenerator8x8[284] = 8'hfe;
assign _c_characterGenerator8x8[285] = 8'h6c;
assign _c_characterGenerator8x8[286] = 8'h6c;
assign _c_characterGenerator8x8[287] = 8'h00;
assign _c_characterGenerator8x8[288] = 8'h30;
assign _c_characterGenerator8x8[289] = 8'h7c;
assign _c_characterGenerator8x8[290] = 8'hc0;
assign _c_characterGenerator8x8[291] = 8'h78;
assign _c_characterGenerator8x8[292] = 8'h0c;
assign _c_characterGenerator8x8[293] = 8'hf8;
assign _c_characterGenerator8x8[294] = 8'h30;
assign _c_characterGenerator8x8[295] = 8'h00;
assign _c_characterGenerator8x8[296] = 8'h00;
assign _c_characterGenerator8x8[297] = 8'hc6;
assign _c_characterGenerator8x8[298] = 8'hcc;
assign _c_characterGenerator8x8[299] = 8'h18;
assign _c_characterGenerator8x8[300] = 8'h30;
assign _c_characterGenerator8x8[301] = 8'h66;
assign _c_characterGenerator8x8[302] = 8'hc6;
assign _c_characterGenerator8x8[303] = 8'h00;
assign _c_characterGenerator8x8[304] = 8'h38;
assign _c_characterGenerator8x8[305] = 8'h6c;
assign _c_characterGenerator8x8[306] = 8'h38;
assign _c_characterGenerator8x8[307] = 8'h76;
assign _c_characterGenerator8x8[308] = 8'hdc;
assign _c_characterGenerator8x8[309] = 8'hcc;
assign _c_characterGenerator8x8[310] = 8'h76;
assign _c_characterGenerator8x8[311] = 8'h00;
assign _c_characterGenerator8x8[312] = 8'h60;
assign _c_characterGenerator8x8[313] = 8'h60;
assign _c_characterGenerator8x8[314] = 8'hc0;
assign _c_characterGenerator8x8[315] = 8'h00;
assign _c_characterGenerator8x8[316] = 8'h00;
assign _c_characterGenerator8x8[317] = 8'h00;
assign _c_characterGenerator8x8[318] = 8'h00;
assign _c_characterGenerator8x8[319] = 8'h00;
assign _c_characterGenerator8x8[320] = 8'h18;
assign _c_characterGenerator8x8[321] = 8'h30;
assign _c_characterGenerator8x8[322] = 8'h60;
assign _c_characterGenerator8x8[323] = 8'h60;
assign _c_characterGenerator8x8[324] = 8'h60;
assign _c_characterGenerator8x8[325] = 8'h30;
assign _c_characterGenerator8x8[326] = 8'h18;
assign _c_characterGenerator8x8[327] = 8'h00;
assign _c_characterGenerator8x8[328] = 8'h60;
assign _c_characterGenerator8x8[329] = 8'h30;
assign _c_characterGenerator8x8[330] = 8'h18;
assign _c_characterGenerator8x8[331] = 8'h18;
assign _c_characterGenerator8x8[332] = 8'h18;
assign _c_characterGenerator8x8[333] = 8'h30;
assign _c_characterGenerator8x8[334] = 8'h60;
assign _c_characterGenerator8x8[335] = 8'h00;
assign _c_characterGenerator8x8[336] = 8'h00;
assign _c_characterGenerator8x8[337] = 8'h66;
assign _c_characterGenerator8x8[338] = 8'h3c;
assign _c_characterGenerator8x8[339] = 8'hff;
assign _c_characterGenerator8x8[340] = 8'h3c;
assign _c_characterGenerator8x8[341] = 8'h66;
assign _c_characterGenerator8x8[342] = 8'h00;
assign _c_characterGenerator8x8[343] = 8'h00;
assign _c_characterGenerator8x8[344] = 8'h00;
assign _c_characterGenerator8x8[345] = 8'h30;
assign _c_characterGenerator8x8[346] = 8'h30;
assign _c_characterGenerator8x8[347] = 8'hfc;
assign _c_characterGenerator8x8[348] = 8'h30;
assign _c_characterGenerator8x8[349] = 8'h30;
assign _c_characterGenerator8x8[350] = 8'h00;
assign _c_characterGenerator8x8[351] = 8'h00;
assign _c_characterGenerator8x8[352] = 8'h00;
assign _c_characterGenerator8x8[353] = 8'h00;
assign _c_characterGenerator8x8[354] = 8'h00;
assign _c_characterGenerator8x8[355] = 8'h00;
assign _c_characterGenerator8x8[356] = 8'h00;
assign _c_characterGenerator8x8[357] = 8'h30;
assign _c_characterGenerator8x8[358] = 8'h30;
assign _c_characterGenerator8x8[359] = 8'h60;
assign _c_characterGenerator8x8[360] = 8'h00;
assign _c_characterGenerator8x8[361] = 8'h00;
assign _c_characterGenerator8x8[362] = 8'h00;
assign _c_characterGenerator8x8[363] = 8'hfc;
assign _c_characterGenerator8x8[364] = 8'h00;
assign _c_characterGenerator8x8[365] = 8'h00;
assign _c_characterGenerator8x8[366] = 8'h00;
assign _c_characterGenerator8x8[367] = 8'h00;
assign _c_characterGenerator8x8[368] = 8'h00;
assign _c_characterGenerator8x8[369] = 8'h00;
assign _c_characterGenerator8x8[370] = 8'h00;
assign _c_characterGenerator8x8[371] = 8'h00;
assign _c_characterGenerator8x8[372] = 8'h00;
assign _c_characterGenerator8x8[373] = 8'h30;
assign _c_characterGenerator8x8[374] = 8'h30;
assign _c_characterGenerator8x8[375] = 8'h00;
assign _c_characterGenerator8x8[376] = 8'h06;
assign _c_characterGenerator8x8[377] = 8'h0c;
assign _c_characterGenerator8x8[378] = 8'h18;
assign _c_characterGenerator8x8[379] = 8'h30;
assign _c_characterGenerator8x8[380] = 8'h60;
assign _c_characterGenerator8x8[381] = 8'hc0;
assign _c_characterGenerator8x8[382] = 8'h80;
assign _c_characterGenerator8x8[383] = 8'h00;
assign _c_characterGenerator8x8[384] = 8'h7c;
assign _c_characterGenerator8x8[385] = 8'hc6;
assign _c_characterGenerator8x8[386] = 8'hce;
assign _c_characterGenerator8x8[387] = 8'hde;
assign _c_characterGenerator8x8[388] = 8'hf6;
assign _c_characterGenerator8x8[389] = 8'he6;
assign _c_characterGenerator8x8[390] = 8'h7c;
assign _c_characterGenerator8x8[391] = 8'h00;
assign _c_characterGenerator8x8[392] = 8'h30;
assign _c_characterGenerator8x8[393] = 8'h70;
assign _c_characterGenerator8x8[394] = 8'h30;
assign _c_characterGenerator8x8[395] = 8'h30;
assign _c_characterGenerator8x8[396] = 8'h30;
assign _c_characterGenerator8x8[397] = 8'h30;
assign _c_characterGenerator8x8[398] = 8'hfc;
assign _c_characterGenerator8x8[399] = 8'h00;
assign _c_characterGenerator8x8[400] = 8'h78;
assign _c_characterGenerator8x8[401] = 8'hcc;
assign _c_characterGenerator8x8[402] = 8'h0c;
assign _c_characterGenerator8x8[403] = 8'h38;
assign _c_characterGenerator8x8[404] = 8'h60;
assign _c_characterGenerator8x8[405] = 8'hcc;
assign _c_characterGenerator8x8[406] = 8'hfc;
assign _c_characterGenerator8x8[407] = 8'h00;
assign _c_characterGenerator8x8[408] = 8'h78;
assign _c_characterGenerator8x8[409] = 8'hcc;
assign _c_characterGenerator8x8[410] = 8'h0c;
assign _c_characterGenerator8x8[411] = 8'h38;
assign _c_characterGenerator8x8[412] = 8'h0c;
assign _c_characterGenerator8x8[413] = 8'hcc;
assign _c_characterGenerator8x8[414] = 8'h78;
assign _c_characterGenerator8x8[415] = 8'h00;
assign _c_characterGenerator8x8[416] = 8'h1c;
assign _c_characterGenerator8x8[417] = 8'h3c;
assign _c_characterGenerator8x8[418] = 8'h6c;
assign _c_characterGenerator8x8[419] = 8'hcc;
assign _c_characterGenerator8x8[420] = 8'hfe;
assign _c_characterGenerator8x8[421] = 8'h0c;
assign _c_characterGenerator8x8[422] = 8'h1e;
assign _c_characterGenerator8x8[423] = 8'h00;
assign _c_characterGenerator8x8[424] = 8'hfc;
assign _c_characterGenerator8x8[425] = 8'hc0;
assign _c_characterGenerator8x8[426] = 8'hf8;
assign _c_characterGenerator8x8[427] = 8'h0c;
assign _c_characterGenerator8x8[428] = 8'h0c;
assign _c_characterGenerator8x8[429] = 8'hcc;
assign _c_characterGenerator8x8[430] = 8'h78;
assign _c_characterGenerator8x8[431] = 8'h00;
assign _c_characterGenerator8x8[432] = 8'h38;
assign _c_characterGenerator8x8[433] = 8'h60;
assign _c_characterGenerator8x8[434] = 8'hc0;
assign _c_characterGenerator8x8[435] = 8'hf8;
assign _c_characterGenerator8x8[436] = 8'hcc;
assign _c_characterGenerator8x8[437] = 8'hcc;
assign _c_characterGenerator8x8[438] = 8'h78;
assign _c_characterGenerator8x8[439] = 8'h00;
assign _c_characterGenerator8x8[440] = 8'hfc;
assign _c_characterGenerator8x8[441] = 8'hcc;
assign _c_characterGenerator8x8[442] = 8'h0c;
assign _c_characterGenerator8x8[443] = 8'h18;
assign _c_characterGenerator8x8[444] = 8'h30;
assign _c_characterGenerator8x8[445] = 8'h30;
assign _c_characterGenerator8x8[446] = 8'h30;
assign _c_characterGenerator8x8[447] = 8'h00;
assign _c_characterGenerator8x8[448] = 8'h78;
assign _c_characterGenerator8x8[449] = 8'hcc;
assign _c_characterGenerator8x8[450] = 8'hcc;
assign _c_characterGenerator8x8[451] = 8'h78;
assign _c_characterGenerator8x8[452] = 8'hcc;
assign _c_characterGenerator8x8[453] = 8'hcc;
assign _c_characterGenerator8x8[454] = 8'h78;
assign _c_characterGenerator8x8[455] = 8'h00;
assign _c_characterGenerator8x8[456] = 8'h78;
assign _c_characterGenerator8x8[457] = 8'hcc;
assign _c_characterGenerator8x8[458] = 8'hcc;
assign _c_characterGenerator8x8[459] = 8'h7c;
assign _c_characterGenerator8x8[460] = 8'h0c;
assign _c_characterGenerator8x8[461] = 8'h18;
assign _c_characterGenerator8x8[462] = 8'h70;
assign _c_characterGenerator8x8[463] = 8'h00;
assign _c_characterGenerator8x8[464] = 8'h00;
assign _c_characterGenerator8x8[465] = 8'h30;
assign _c_characterGenerator8x8[466] = 8'h30;
assign _c_characterGenerator8x8[467] = 8'h00;
assign _c_characterGenerator8x8[468] = 8'h00;
assign _c_characterGenerator8x8[469] = 8'h30;
assign _c_characterGenerator8x8[470] = 8'h30;
assign _c_characterGenerator8x8[471] = 8'h00;
assign _c_characterGenerator8x8[472] = 8'h00;
assign _c_characterGenerator8x8[473] = 8'h30;
assign _c_characterGenerator8x8[474] = 8'h30;
assign _c_characterGenerator8x8[475] = 8'h00;
assign _c_characterGenerator8x8[476] = 8'h00;
assign _c_characterGenerator8x8[477] = 8'h30;
assign _c_characterGenerator8x8[478] = 8'h30;
assign _c_characterGenerator8x8[479] = 8'h60;
assign _c_characterGenerator8x8[480] = 8'h18;
assign _c_characterGenerator8x8[481] = 8'h30;
assign _c_characterGenerator8x8[482] = 8'h60;
assign _c_characterGenerator8x8[483] = 8'hc0;
assign _c_characterGenerator8x8[484] = 8'h60;
assign _c_characterGenerator8x8[485] = 8'h30;
assign _c_characterGenerator8x8[486] = 8'h18;
assign _c_characterGenerator8x8[487] = 8'h00;
assign _c_characterGenerator8x8[488] = 8'h00;
assign _c_characterGenerator8x8[489] = 8'h00;
assign _c_characterGenerator8x8[490] = 8'hfc;
assign _c_characterGenerator8x8[491] = 8'h00;
assign _c_characterGenerator8x8[492] = 8'h00;
assign _c_characterGenerator8x8[493] = 8'hfc;
assign _c_characterGenerator8x8[494] = 8'h00;
assign _c_characterGenerator8x8[495] = 8'h00;
assign _c_characterGenerator8x8[496] = 8'h60;
assign _c_characterGenerator8x8[497] = 8'h30;
assign _c_characterGenerator8x8[498] = 8'h18;
assign _c_characterGenerator8x8[499] = 8'h0c;
assign _c_characterGenerator8x8[500] = 8'h18;
assign _c_characterGenerator8x8[501] = 8'h30;
assign _c_characterGenerator8x8[502] = 8'h60;
assign _c_characterGenerator8x8[503] = 8'h00;
assign _c_characterGenerator8x8[504] = 8'h78;
assign _c_characterGenerator8x8[505] = 8'hcc;
assign _c_characterGenerator8x8[506] = 8'h0c;
assign _c_characterGenerator8x8[507] = 8'h18;
assign _c_characterGenerator8x8[508] = 8'h30;
assign _c_characterGenerator8x8[509] = 8'h00;
assign _c_characterGenerator8x8[510] = 8'h30;
assign _c_characterGenerator8x8[511] = 8'h00;
assign _c_characterGenerator8x8[512] = 8'h7c;
assign _c_characterGenerator8x8[513] = 8'hc6;
assign _c_characterGenerator8x8[514] = 8'hde;
assign _c_characterGenerator8x8[515] = 8'hde;
assign _c_characterGenerator8x8[516] = 8'hde;
assign _c_characterGenerator8x8[517] = 8'hc0;
assign _c_characterGenerator8x8[518] = 8'h78;
assign _c_characterGenerator8x8[519] = 8'h00;
assign _c_characterGenerator8x8[520] = 8'h30;
assign _c_characterGenerator8x8[521] = 8'h78;
assign _c_characterGenerator8x8[522] = 8'hcc;
assign _c_characterGenerator8x8[523] = 8'hcc;
assign _c_characterGenerator8x8[524] = 8'hfc;
assign _c_characterGenerator8x8[525] = 8'hcc;
assign _c_characterGenerator8x8[526] = 8'hcc;
assign _c_characterGenerator8x8[527] = 8'h00;
assign _c_characterGenerator8x8[528] = 8'hfc;
assign _c_characterGenerator8x8[529] = 8'h66;
assign _c_characterGenerator8x8[530] = 8'h66;
assign _c_characterGenerator8x8[531] = 8'h7c;
assign _c_characterGenerator8x8[532] = 8'h66;
assign _c_characterGenerator8x8[533] = 8'h66;
assign _c_characterGenerator8x8[534] = 8'hfc;
assign _c_characterGenerator8x8[535] = 8'h00;
assign _c_characterGenerator8x8[536] = 8'h3c;
assign _c_characterGenerator8x8[537] = 8'h66;
assign _c_characterGenerator8x8[538] = 8'hc0;
assign _c_characterGenerator8x8[539] = 8'hc0;
assign _c_characterGenerator8x8[540] = 8'hc0;
assign _c_characterGenerator8x8[541] = 8'h66;
assign _c_characterGenerator8x8[542] = 8'h3c;
assign _c_characterGenerator8x8[543] = 8'h00;
assign _c_characterGenerator8x8[544] = 8'hf8;
assign _c_characterGenerator8x8[545] = 8'h6c;
assign _c_characterGenerator8x8[546] = 8'h66;
assign _c_characterGenerator8x8[547] = 8'h66;
assign _c_characterGenerator8x8[548] = 8'h66;
assign _c_characterGenerator8x8[549] = 8'h6c;
assign _c_characterGenerator8x8[550] = 8'hf8;
assign _c_characterGenerator8x8[551] = 8'h00;
assign _c_characterGenerator8x8[552] = 8'hfe;
assign _c_characterGenerator8x8[553] = 8'h62;
assign _c_characterGenerator8x8[554] = 8'h68;
assign _c_characterGenerator8x8[555] = 8'h78;
assign _c_characterGenerator8x8[556] = 8'h68;
assign _c_characterGenerator8x8[557] = 8'h62;
assign _c_characterGenerator8x8[558] = 8'hfe;
assign _c_characterGenerator8x8[559] = 8'h00;
assign _c_characterGenerator8x8[560] = 8'hfe;
assign _c_characterGenerator8x8[561] = 8'h62;
assign _c_characterGenerator8x8[562] = 8'h68;
assign _c_characterGenerator8x8[563] = 8'h78;
assign _c_characterGenerator8x8[564] = 8'h68;
assign _c_characterGenerator8x8[565] = 8'h60;
assign _c_characterGenerator8x8[566] = 8'hf0;
assign _c_characterGenerator8x8[567] = 8'h00;
assign _c_characterGenerator8x8[568] = 8'h3c;
assign _c_characterGenerator8x8[569] = 8'h66;
assign _c_characterGenerator8x8[570] = 8'hc0;
assign _c_characterGenerator8x8[571] = 8'hc0;
assign _c_characterGenerator8x8[572] = 8'hce;
assign _c_characterGenerator8x8[573] = 8'h66;
assign _c_characterGenerator8x8[574] = 8'h3e;
assign _c_characterGenerator8x8[575] = 8'h00;
assign _c_characterGenerator8x8[576] = 8'hcc;
assign _c_characterGenerator8x8[577] = 8'hcc;
assign _c_characterGenerator8x8[578] = 8'hcc;
assign _c_characterGenerator8x8[579] = 8'hfc;
assign _c_characterGenerator8x8[580] = 8'hcc;
assign _c_characterGenerator8x8[581] = 8'hcc;
assign _c_characterGenerator8x8[582] = 8'hcc;
assign _c_characterGenerator8x8[583] = 8'h00;
assign _c_characterGenerator8x8[584] = 8'h78;
assign _c_characterGenerator8x8[585] = 8'h30;
assign _c_characterGenerator8x8[586] = 8'h30;
assign _c_characterGenerator8x8[587] = 8'h30;
assign _c_characterGenerator8x8[588] = 8'h30;
assign _c_characterGenerator8x8[589] = 8'h30;
assign _c_characterGenerator8x8[590] = 8'h78;
assign _c_characterGenerator8x8[591] = 8'h00;
assign _c_characterGenerator8x8[592] = 8'h1e;
assign _c_characterGenerator8x8[593] = 8'h0c;
assign _c_characterGenerator8x8[594] = 8'h0c;
assign _c_characterGenerator8x8[595] = 8'h0c;
assign _c_characterGenerator8x8[596] = 8'hcc;
assign _c_characterGenerator8x8[597] = 8'hcc;
assign _c_characterGenerator8x8[598] = 8'h78;
assign _c_characterGenerator8x8[599] = 8'h00;
assign _c_characterGenerator8x8[600] = 8'he6;
assign _c_characterGenerator8x8[601] = 8'h66;
assign _c_characterGenerator8x8[602] = 8'h6c;
assign _c_characterGenerator8x8[603] = 8'h78;
assign _c_characterGenerator8x8[604] = 8'h6c;
assign _c_characterGenerator8x8[605] = 8'h66;
assign _c_characterGenerator8x8[606] = 8'he6;
assign _c_characterGenerator8x8[607] = 8'h00;
assign _c_characterGenerator8x8[608] = 8'hf0;
assign _c_characterGenerator8x8[609] = 8'h60;
assign _c_characterGenerator8x8[610] = 8'h60;
assign _c_characterGenerator8x8[611] = 8'h60;
assign _c_characterGenerator8x8[612] = 8'h62;
assign _c_characterGenerator8x8[613] = 8'h66;
assign _c_characterGenerator8x8[614] = 8'hfe;
assign _c_characterGenerator8x8[615] = 8'h00;
assign _c_characterGenerator8x8[616] = 8'hc6;
assign _c_characterGenerator8x8[617] = 8'hee;
assign _c_characterGenerator8x8[618] = 8'hfe;
assign _c_characterGenerator8x8[619] = 8'hfe;
assign _c_characterGenerator8x8[620] = 8'hd6;
assign _c_characterGenerator8x8[621] = 8'hc6;
assign _c_characterGenerator8x8[622] = 8'hc6;
assign _c_characterGenerator8x8[623] = 8'h00;
assign _c_characterGenerator8x8[624] = 8'hc6;
assign _c_characterGenerator8x8[625] = 8'he6;
assign _c_characterGenerator8x8[626] = 8'hf6;
assign _c_characterGenerator8x8[627] = 8'hde;
assign _c_characterGenerator8x8[628] = 8'hce;
assign _c_characterGenerator8x8[629] = 8'hc6;
assign _c_characterGenerator8x8[630] = 8'hc6;
assign _c_characterGenerator8x8[631] = 8'h00;
assign _c_characterGenerator8x8[632] = 8'h38;
assign _c_characterGenerator8x8[633] = 8'h6c;
assign _c_characterGenerator8x8[634] = 8'hc6;
assign _c_characterGenerator8x8[635] = 8'hc6;
assign _c_characterGenerator8x8[636] = 8'hc6;
assign _c_characterGenerator8x8[637] = 8'h6c;
assign _c_characterGenerator8x8[638] = 8'h38;
assign _c_characterGenerator8x8[639] = 8'h00;
assign _c_characterGenerator8x8[640] = 8'hfc;
assign _c_characterGenerator8x8[641] = 8'h66;
assign _c_characterGenerator8x8[642] = 8'h66;
assign _c_characterGenerator8x8[643] = 8'h7c;
assign _c_characterGenerator8x8[644] = 8'h60;
assign _c_characterGenerator8x8[645] = 8'h60;
assign _c_characterGenerator8x8[646] = 8'hf0;
assign _c_characterGenerator8x8[647] = 8'h00;
assign _c_characterGenerator8x8[648] = 8'h78;
assign _c_characterGenerator8x8[649] = 8'hcc;
assign _c_characterGenerator8x8[650] = 8'hcc;
assign _c_characterGenerator8x8[651] = 8'hcc;
assign _c_characterGenerator8x8[652] = 8'hdc;
assign _c_characterGenerator8x8[653] = 8'h78;
assign _c_characterGenerator8x8[654] = 8'h1c;
assign _c_characterGenerator8x8[655] = 8'h00;
assign _c_characterGenerator8x8[656] = 8'hfc;
assign _c_characterGenerator8x8[657] = 8'h66;
assign _c_characterGenerator8x8[658] = 8'h66;
assign _c_characterGenerator8x8[659] = 8'h7c;
assign _c_characterGenerator8x8[660] = 8'h6c;
assign _c_characterGenerator8x8[661] = 8'h66;
assign _c_characterGenerator8x8[662] = 8'he6;
assign _c_characterGenerator8x8[663] = 8'h00;
assign _c_characterGenerator8x8[664] = 8'h78;
assign _c_characterGenerator8x8[665] = 8'hcc;
assign _c_characterGenerator8x8[666] = 8'he0;
assign _c_characterGenerator8x8[667] = 8'h70;
assign _c_characterGenerator8x8[668] = 8'h1c;
assign _c_characterGenerator8x8[669] = 8'hcc;
assign _c_characterGenerator8x8[670] = 8'h78;
assign _c_characterGenerator8x8[671] = 8'h00;
assign _c_characterGenerator8x8[672] = 8'hfc;
assign _c_characterGenerator8x8[673] = 8'hb4;
assign _c_characterGenerator8x8[674] = 8'h30;
assign _c_characterGenerator8x8[675] = 8'h30;
assign _c_characterGenerator8x8[676] = 8'h30;
assign _c_characterGenerator8x8[677] = 8'h30;
assign _c_characterGenerator8x8[678] = 8'h78;
assign _c_characterGenerator8x8[679] = 8'h00;
assign _c_characterGenerator8x8[680] = 8'hcc;
assign _c_characterGenerator8x8[681] = 8'hcc;
assign _c_characterGenerator8x8[682] = 8'hcc;
assign _c_characterGenerator8x8[683] = 8'hcc;
assign _c_characterGenerator8x8[684] = 8'hcc;
assign _c_characterGenerator8x8[685] = 8'hcc;
assign _c_characterGenerator8x8[686] = 8'hfc;
assign _c_characterGenerator8x8[687] = 8'h00;
assign _c_characterGenerator8x8[688] = 8'hcc;
assign _c_characterGenerator8x8[689] = 8'hcc;
assign _c_characterGenerator8x8[690] = 8'hcc;
assign _c_characterGenerator8x8[691] = 8'hcc;
assign _c_characterGenerator8x8[692] = 8'hcc;
assign _c_characterGenerator8x8[693] = 8'h78;
assign _c_characterGenerator8x8[694] = 8'h30;
assign _c_characterGenerator8x8[695] = 8'h00;
assign _c_characterGenerator8x8[696] = 8'hc6;
assign _c_characterGenerator8x8[697] = 8'hc6;
assign _c_characterGenerator8x8[698] = 8'hc6;
assign _c_characterGenerator8x8[699] = 8'hd6;
assign _c_characterGenerator8x8[700] = 8'hfe;
assign _c_characterGenerator8x8[701] = 8'hee;
assign _c_characterGenerator8x8[702] = 8'hc6;
assign _c_characterGenerator8x8[703] = 8'h00;
assign _c_characterGenerator8x8[704] = 8'hc6;
assign _c_characterGenerator8x8[705] = 8'hc6;
assign _c_characterGenerator8x8[706] = 8'h6c;
assign _c_characterGenerator8x8[707] = 8'h38;
assign _c_characterGenerator8x8[708] = 8'h38;
assign _c_characterGenerator8x8[709] = 8'h6c;
assign _c_characterGenerator8x8[710] = 8'hc6;
assign _c_characterGenerator8x8[711] = 8'h00;
assign _c_characterGenerator8x8[712] = 8'hcc;
assign _c_characterGenerator8x8[713] = 8'hcc;
assign _c_characterGenerator8x8[714] = 8'hcc;
assign _c_characterGenerator8x8[715] = 8'h78;
assign _c_characterGenerator8x8[716] = 8'h30;
assign _c_characterGenerator8x8[717] = 8'h30;
assign _c_characterGenerator8x8[718] = 8'h78;
assign _c_characterGenerator8x8[719] = 8'h00;
assign _c_characterGenerator8x8[720] = 8'hfe;
assign _c_characterGenerator8x8[721] = 8'hc6;
assign _c_characterGenerator8x8[722] = 8'h8c;
assign _c_characterGenerator8x8[723] = 8'h18;
assign _c_characterGenerator8x8[724] = 8'h32;
assign _c_characterGenerator8x8[725] = 8'h66;
assign _c_characterGenerator8x8[726] = 8'hfe;
assign _c_characterGenerator8x8[727] = 8'h00;
assign _c_characterGenerator8x8[728] = 8'h78;
assign _c_characterGenerator8x8[729] = 8'h60;
assign _c_characterGenerator8x8[730] = 8'h60;
assign _c_characterGenerator8x8[731] = 8'h60;
assign _c_characterGenerator8x8[732] = 8'h60;
assign _c_characterGenerator8x8[733] = 8'h60;
assign _c_characterGenerator8x8[734] = 8'h78;
assign _c_characterGenerator8x8[735] = 8'h00;
assign _c_characterGenerator8x8[736] = 8'hc0;
assign _c_characterGenerator8x8[737] = 8'h60;
assign _c_characterGenerator8x8[738] = 8'h30;
assign _c_characterGenerator8x8[739] = 8'h18;
assign _c_characterGenerator8x8[740] = 8'h0c;
assign _c_characterGenerator8x8[741] = 8'h06;
assign _c_characterGenerator8x8[742] = 8'h02;
assign _c_characterGenerator8x8[743] = 8'h00;
assign _c_characterGenerator8x8[744] = 8'h78;
assign _c_characterGenerator8x8[745] = 8'h18;
assign _c_characterGenerator8x8[746] = 8'h18;
assign _c_characterGenerator8x8[747] = 8'h18;
assign _c_characterGenerator8x8[748] = 8'h18;
assign _c_characterGenerator8x8[749] = 8'h18;
assign _c_characterGenerator8x8[750] = 8'h78;
assign _c_characterGenerator8x8[751] = 8'h00;
assign _c_characterGenerator8x8[752] = 8'h10;
assign _c_characterGenerator8x8[753] = 8'h38;
assign _c_characterGenerator8x8[754] = 8'h6c;
assign _c_characterGenerator8x8[755] = 8'hc6;
assign _c_characterGenerator8x8[756] = 8'h00;
assign _c_characterGenerator8x8[757] = 8'h00;
assign _c_characterGenerator8x8[758] = 8'h00;
assign _c_characterGenerator8x8[759] = 8'h00;
assign _c_characterGenerator8x8[760] = 8'h00;
assign _c_characterGenerator8x8[761] = 8'h00;
assign _c_characterGenerator8x8[762] = 8'h00;
assign _c_characterGenerator8x8[763] = 8'h00;
assign _c_characterGenerator8x8[764] = 8'h00;
assign _c_characterGenerator8x8[765] = 8'h00;
assign _c_characterGenerator8x8[766] = 8'h00;
assign _c_characterGenerator8x8[767] = 8'hff;
assign _c_characterGenerator8x8[768] = 8'h30;
assign _c_characterGenerator8x8[769] = 8'h30;
assign _c_characterGenerator8x8[770] = 8'h18;
assign _c_characterGenerator8x8[771] = 8'h00;
assign _c_characterGenerator8x8[772] = 8'h00;
assign _c_characterGenerator8x8[773] = 8'h00;
assign _c_characterGenerator8x8[774] = 8'h00;
assign _c_characterGenerator8x8[775] = 8'h00;
assign _c_characterGenerator8x8[776] = 8'h00;
assign _c_characterGenerator8x8[777] = 8'h00;
assign _c_characterGenerator8x8[778] = 8'h78;
assign _c_characterGenerator8x8[779] = 8'h0c;
assign _c_characterGenerator8x8[780] = 8'h7c;
assign _c_characterGenerator8x8[781] = 8'hcc;
assign _c_characterGenerator8x8[782] = 8'h76;
assign _c_characterGenerator8x8[783] = 8'h00;
assign _c_characterGenerator8x8[784] = 8'he0;
assign _c_characterGenerator8x8[785] = 8'h60;
assign _c_characterGenerator8x8[786] = 8'h60;
assign _c_characterGenerator8x8[787] = 8'h7c;
assign _c_characterGenerator8x8[788] = 8'h66;
assign _c_characterGenerator8x8[789] = 8'h66;
assign _c_characterGenerator8x8[790] = 8'hdc;
assign _c_characterGenerator8x8[791] = 8'h00;
assign _c_characterGenerator8x8[792] = 8'h00;
assign _c_characterGenerator8x8[793] = 8'h00;
assign _c_characterGenerator8x8[794] = 8'h78;
assign _c_characterGenerator8x8[795] = 8'hcc;
assign _c_characterGenerator8x8[796] = 8'hc0;
assign _c_characterGenerator8x8[797] = 8'hcc;
assign _c_characterGenerator8x8[798] = 8'h78;
assign _c_characterGenerator8x8[799] = 8'h00;
assign _c_characterGenerator8x8[800] = 8'h1c;
assign _c_characterGenerator8x8[801] = 8'h0c;
assign _c_characterGenerator8x8[802] = 8'h0c;
assign _c_characterGenerator8x8[803] = 8'h7c;
assign _c_characterGenerator8x8[804] = 8'hcc;
assign _c_characterGenerator8x8[805] = 8'hcc;
assign _c_characterGenerator8x8[806] = 8'h76;
assign _c_characterGenerator8x8[807] = 8'h00;
assign _c_characterGenerator8x8[808] = 8'h00;
assign _c_characterGenerator8x8[809] = 8'h00;
assign _c_characterGenerator8x8[810] = 8'h78;
assign _c_characterGenerator8x8[811] = 8'hcc;
assign _c_characterGenerator8x8[812] = 8'hfc;
assign _c_characterGenerator8x8[813] = 8'hc0;
assign _c_characterGenerator8x8[814] = 8'h78;
assign _c_characterGenerator8x8[815] = 8'h00;
assign _c_characterGenerator8x8[816] = 8'h38;
assign _c_characterGenerator8x8[817] = 8'h6c;
assign _c_characterGenerator8x8[818] = 8'h60;
assign _c_characterGenerator8x8[819] = 8'hf0;
assign _c_characterGenerator8x8[820] = 8'h60;
assign _c_characterGenerator8x8[821] = 8'h60;
assign _c_characterGenerator8x8[822] = 8'hf0;
assign _c_characterGenerator8x8[823] = 8'h00;
assign _c_characterGenerator8x8[824] = 8'h00;
assign _c_characterGenerator8x8[825] = 8'h00;
assign _c_characterGenerator8x8[826] = 8'h76;
assign _c_characterGenerator8x8[827] = 8'hcc;
assign _c_characterGenerator8x8[828] = 8'hcc;
assign _c_characterGenerator8x8[829] = 8'h7c;
assign _c_characterGenerator8x8[830] = 8'h0c;
assign _c_characterGenerator8x8[831] = 8'hf8;
assign _c_characterGenerator8x8[832] = 8'he0;
assign _c_characterGenerator8x8[833] = 8'h60;
assign _c_characterGenerator8x8[834] = 8'h6c;
assign _c_characterGenerator8x8[835] = 8'h76;
assign _c_characterGenerator8x8[836] = 8'h66;
assign _c_characterGenerator8x8[837] = 8'h66;
assign _c_characterGenerator8x8[838] = 8'he6;
assign _c_characterGenerator8x8[839] = 8'h00;
assign _c_characterGenerator8x8[840] = 8'h30;
assign _c_characterGenerator8x8[841] = 8'h00;
assign _c_characterGenerator8x8[842] = 8'h70;
assign _c_characterGenerator8x8[843] = 8'h30;
assign _c_characterGenerator8x8[844] = 8'h30;
assign _c_characterGenerator8x8[845] = 8'h30;
assign _c_characterGenerator8x8[846] = 8'h78;
assign _c_characterGenerator8x8[847] = 8'h00;
assign _c_characterGenerator8x8[848] = 8'h0c;
assign _c_characterGenerator8x8[849] = 8'h00;
assign _c_characterGenerator8x8[850] = 8'h0c;
assign _c_characterGenerator8x8[851] = 8'h0c;
assign _c_characterGenerator8x8[852] = 8'h0c;
assign _c_characterGenerator8x8[853] = 8'hcc;
assign _c_characterGenerator8x8[854] = 8'hcc;
assign _c_characterGenerator8x8[855] = 8'h78;
assign _c_characterGenerator8x8[856] = 8'he0;
assign _c_characterGenerator8x8[857] = 8'h60;
assign _c_characterGenerator8x8[858] = 8'h66;
assign _c_characterGenerator8x8[859] = 8'h6c;
assign _c_characterGenerator8x8[860] = 8'h78;
assign _c_characterGenerator8x8[861] = 8'h6c;
assign _c_characterGenerator8x8[862] = 8'he6;
assign _c_characterGenerator8x8[863] = 8'h00;
assign _c_characterGenerator8x8[864] = 8'h70;
assign _c_characterGenerator8x8[865] = 8'h30;
assign _c_characterGenerator8x8[866] = 8'h30;
assign _c_characterGenerator8x8[867] = 8'h30;
assign _c_characterGenerator8x8[868] = 8'h30;
assign _c_characterGenerator8x8[869] = 8'h30;
assign _c_characterGenerator8x8[870] = 8'h78;
assign _c_characterGenerator8x8[871] = 8'h00;
assign _c_characterGenerator8x8[872] = 8'h00;
assign _c_characterGenerator8x8[873] = 8'h00;
assign _c_characterGenerator8x8[874] = 8'hcc;
assign _c_characterGenerator8x8[875] = 8'hfe;
assign _c_characterGenerator8x8[876] = 8'hfe;
assign _c_characterGenerator8x8[877] = 8'hd6;
assign _c_characterGenerator8x8[878] = 8'hc6;
assign _c_characterGenerator8x8[879] = 8'h00;
assign _c_characterGenerator8x8[880] = 8'h00;
assign _c_characterGenerator8x8[881] = 8'h00;
assign _c_characterGenerator8x8[882] = 8'hf8;
assign _c_characterGenerator8x8[883] = 8'hcc;
assign _c_characterGenerator8x8[884] = 8'hcc;
assign _c_characterGenerator8x8[885] = 8'hcc;
assign _c_characterGenerator8x8[886] = 8'hcc;
assign _c_characterGenerator8x8[887] = 8'h00;
assign _c_characterGenerator8x8[888] = 8'h00;
assign _c_characterGenerator8x8[889] = 8'h00;
assign _c_characterGenerator8x8[890] = 8'h78;
assign _c_characterGenerator8x8[891] = 8'hcc;
assign _c_characterGenerator8x8[892] = 8'hcc;
assign _c_characterGenerator8x8[893] = 8'hcc;
assign _c_characterGenerator8x8[894] = 8'h78;
assign _c_characterGenerator8x8[895] = 8'h00;
assign _c_characterGenerator8x8[896] = 8'h00;
assign _c_characterGenerator8x8[897] = 8'h00;
assign _c_characterGenerator8x8[898] = 8'hdc;
assign _c_characterGenerator8x8[899] = 8'h66;
assign _c_characterGenerator8x8[900] = 8'h66;
assign _c_characterGenerator8x8[901] = 8'h7c;
assign _c_characterGenerator8x8[902] = 8'h60;
assign _c_characterGenerator8x8[903] = 8'hf0;
assign _c_characterGenerator8x8[904] = 8'h00;
assign _c_characterGenerator8x8[905] = 8'h00;
assign _c_characterGenerator8x8[906] = 8'h76;
assign _c_characterGenerator8x8[907] = 8'hcc;
assign _c_characterGenerator8x8[908] = 8'hcc;
assign _c_characterGenerator8x8[909] = 8'h7c;
assign _c_characterGenerator8x8[910] = 8'h0c;
assign _c_characterGenerator8x8[911] = 8'h1e;
assign _c_characterGenerator8x8[912] = 8'h00;
assign _c_characterGenerator8x8[913] = 8'h00;
assign _c_characterGenerator8x8[914] = 8'hdc;
assign _c_characterGenerator8x8[915] = 8'h76;
assign _c_characterGenerator8x8[916] = 8'h66;
assign _c_characterGenerator8x8[917] = 8'h60;
assign _c_characterGenerator8x8[918] = 8'hf0;
assign _c_characterGenerator8x8[919] = 8'h00;
assign _c_characterGenerator8x8[920] = 8'h00;
assign _c_characterGenerator8x8[921] = 8'h00;
assign _c_characterGenerator8x8[922] = 8'h7c;
assign _c_characterGenerator8x8[923] = 8'hc0;
assign _c_characterGenerator8x8[924] = 8'h78;
assign _c_characterGenerator8x8[925] = 8'h0c;
assign _c_characterGenerator8x8[926] = 8'hf8;
assign _c_characterGenerator8x8[927] = 8'h00;
assign _c_characterGenerator8x8[928] = 8'h10;
assign _c_characterGenerator8x8[929] = 8'h30;
assign _c_characterGenerator8x8[930] = 8'h7c;
assign _c_characterGenerator8x8[931] = 8'h30;
assign _c_characterGenerator8x8[932] = 8'h30;
assign _c_characterGenerator8x8[933] = 8'h34;
assign _c_characterGenerator8x8[934] = 8'h18;
assign _c_characterGenerator8x8[935] = 8'h00;
assign _c_characterGenerator8x8[936] = 8'h00;
assign _c_characterGenerator8x8[937] = 8'h00;
assign _c_characterGenerator8x8[938] = 8'hcc;
assign _c_characterGenerator8x8[939] = 8'hcc;
assign _c_characterGenerator8x8[940] = 8'hcc;
assign _c_characterGenerator8x8[941] = 8'hcc;
assign _c_characterGenerator8x8[942] = 8'h76;
assign _c_characterGenerator8x8[943] = 8'h00;
assign _c_characterGenerator8x8[944] = 8'h00;
assign _c_characterGenerator8x8[945] = 8'h00;
assign _c_characterGenerator8x8[946] = 8'hcc;
assign _c_characterGenerator8x8[947] = 8'hcc;
assign _c_characterGenerator8x8[948] = 8'hcc;
assign _c_characterGenerator8x8[949] = 8'h78;
assign _c_characterGenerator8x8[950] = 8'h30;
assign _c_characterGenerator8x8[951] = 8'h00;
assign _c_characterGenerator8x8[952] = 8'h00;
assign _c_characterGenerator8x8[953] = 8'h00;
assign _c_characterGenerator8x8[954] = 8'hc6;
assign _c_characterGenerator8x8[955] = 8'hd6;
assign _c_characterGenerator8x8[956] = 8'hfe;
assign _c_characterGenerator8x8[957] = 8'hfe;
assign _c_characterGenerator8x8[958] = 8'h6c;
assign _c_characterGenerator8x8[959] = 8'h00;
assign _c_characterGenerator8x8[960] = 8'h00;
assign _c_characterGenerator8x8[961] = 8'h00;
assign _c_characterGenerator8x8[962] = 8'hc6;
assign _c_characterGenerator8x8[963] = 8'h6c;
assign _c_characterGenerator8x8[964] = 8'h38;
assign _c_characterGenerator8x8[965] = 8'h6c;
assign _c_characterGenerator8x8[966] = 8'hc6;
assign _c_characterGenerator8x8[967] = 8'h00;
assign _c_characterGenerator8x8[968] = 8'h00;
assign _c_characterGenerator8x8[969] = 8'h00;
assign _c_characterGenerator8x8[970] = 8'hcc;
assign _c_characterGenerator8x8[971] = 8'hcc;
assign _c_characterGenerator8x8[972] = 8'hcc;
assign _c_characterGenerator8x8[973] = 8'h7c;
assign _c_characterGenerator8x8[974] = 8'h0c;
assign _c_characterGenerator8x8[975] = 8'hf8;
assign _c_characterGenerator8x8[976] = 8'h00;
assign _c_characterGenerator8x8[977] = 8'h00;
assign _c_characterGenerator8x8[978] = 8'hfc;
assign _c_characterGenerator8x8[979] = 8'h98;
assign _c_characterGenerator8x8[980] = 8'h30;
assign _c_characterGenerator8x8[981] = 8'h64;
assign _c_characterGenerator8x8[982] = 8'hfc;
assign _c_characterGenerator8x8[983] = 8'h00;
assign _c_characterGenerator8x8[984] = 8'h1c;
assign _c_characterGenerator8x8[985] = 8'h30;
assign _c_characterGenerator8x8[986] = 8'h30;
assign _c_characterGenerator8x8[987] = 8'he0;
assign _c_characterGenerator8x8[988] = 8'h30;
assign _c_characterGenerator8x8[989] = 8'h30;
assign _c_characterGenerator8x8[990] = 8'h1c;
assign _c_characterGenerator8x8[991] = 8'h00;
assign _c_characterGenerator8x8[992] = 8'h18;
assign _c_characterGenerator8x8[993] = 8'h18;
assign _c_characterGenerator8x8[994] = 8'h18;
assign _c_characterGenerator8x8[995] = 8'h00;
assign _c_characterGenerator8x8[996] = 8'h18;
assign _c_characterGenerator8x8[997] = 8'h18;
assign _c_characterGenerator8x8[998] = 8'h18;
assign _c_characterGenerator8x8[999] = 8'h00;
assign _c_characterGenerator8x8[1000] = 8'he0;
assign _c_characterGenerator8x8[1001] = 8'h30;
assign _c_characterGenerator8x8[1002] = 8'h30;
assign _c_characterGenerator8x8[1003] = 8'h1c;
assign _c_characterGenerator8x8[1004] = 8'h30;
assign _c_characterGenerator8x8[1005] = 8'h30;
assign _c_characterGenerator8x8[1006] = 8'he0;
assign _c_characterGenerator8x8[1007] = 8'h00;
assign _c_characterGenerator8x8[1008] = 8'h76;
assign _c_characterGenerator8x8[1009] = 8'hdc;
assign _c_characterGenerator8x8[1010] = 8'h00;
assign _c_characterGenerator8x8[1011] = 8'h00;
assign _c_characterGenerator8x8[1012] = 8'h00;
assign _c_characterGenerator8x8[1013] = 8'h00;
assign _c_characterGenerator8x8[1014] = 8'h00;
assign _c_characterGenerator8x8[1015] = 8'h00;
assign _c_characterGenerator8x8[1016] = 8'h00;
assign _c_characterGenerator8x8[1017] = 8'h10;
assign _c_characterGenerator8x8[1018] = 8'h38;
assign _c_characterGenerator8x8[1019] = 8'h6c;
assign _c_characterGenerator8x8[1020] = 8'hc6;
assign _c_characterGenerator8x8[1021] = 8'hc6;
assign _c_characterGenerator8x8[1022] = 8'hfe;
assign _c_characterGenerator8x8[1023] = 8'h00;
assign _c_characterGenerator8x8[1024] = 8'h78;
assign _c_characterGenerator8x8[1025] = 8'hcc;
assign _c_characterGenerator8x8[1026] = 8'hc0;
assign _c_characterGenerator8x8[1027] = 8'hcc;
assign _c_characterGenerator8x8[1028] = 8'h78;
assign _c_characterGenerator8x8[1029] = 8'h18;
assign _c_characterGenerator8x8[1030] = 8'h0c;
assign _c_characterGenerator8x8[1031] = 8'h78;
assign _c_characterGenerator8x8[1032] = 8'h00;
assign _c_characterGenerator8x8[1033] = 8'hcc;
assign _c_characterGenerator8x8[1034] = 8'h00;
assign _c_characterGenerator8x8[1035] = 8'hcc;
assign _c_characterGenerator8x8[1036] = 8'hcc;
assign _c_characterGenerator8x8[1037] = 8'hcc;
assign _c_characterGenerator8x8[1038] = 8'h7e;
assign _c_characterGenerator8x8[1039] = 8'h00;
assign _c_characterGenerator8x8[1040] = 8'h1c;
assign _c_characterGenerator8x8[1041] = 8'h00;
assign _c_characterGenerator8x8[1042] = 8'h78;
assign _c_characterGenerator8x8[1043] = 8'hcc;
assign _c_characterGenerator8x8[1044] = 8'hfc;
assign _c_characterGenerator8x8[1045] = 8'hc0;
assign _c_characterGenerator8x8[1046] = 8'h78;
assign _c_characterGenerator8x8[1047] = 8'h00;
assign _c_characterGenerator8x8[1048] = 8'h7e;
assign _c_characterGenerator8x8[1049] = 8'hc3;
assign _c_characterGenerator8x8[1050] = 8'h3c;
assign _c_characterGenerator8x8[1051] = 8'h06;
assign _c_characterGenerator8x8[1052] = 8'h3e;
assign _c_characterGenerator8x8[1053] = 8'h66;
assign _c_characterGenerator8x8[1054] = 8'h3f;
assign _c_characterGenerator8x8[1055] = 8'h00;
assign _c_characterGenerator8x8[1056] = 8'hcc;
assign _c_characterGenerator8x8[1057] = 8'h00;
assign _c_characterGenerator8x8[1058] = 8'h78;
assign _c_characterGenerator8x8[1059] = 8'h0c;
assign _c_characterGenerator8x8[1060] = 8'h7c;
assign _c_characterGenerator8x8[1061] = 8'hcc;
assign _c_characterGenerator8x8[1062] = 8'h7e;
assign _c_characterGenerator8x8[1063] = 8'h00;
assign _c_characterGenerator8x8[1064] = 8'he0;
assign _c_characterGenerator8x8[1065] = 8'h00;
assign _c_characterGenerator8x8[1066] = 8'h78;
assign _c_characterGenerator8x8[1067] = 8'h0c;
assign _c_characterGenerator8x8[1068] = 8'h7c;
assign _c_characterGenerator8x8[1069] = 8'hcc;
assign _c_characterGenerator8x8[1070] = 8'h7e;
assign _c_characterGenerator8x8[1071] = 8'h00;
assign _c_characterGenerator8x8[1072] = 8'h30;
assign _c_characterGenerator8x8[1073] = 8'h30;
assign _c_characterGenerator8x8[1074] = 8'h78;
assign _c_characterGenerator8x8[1075] = 8'h0c;
assign _c_characterGenerator8x8[1076] = 8'h7c;
assign _c_characterGenerator8x8[1077] = 8'hcc;
assign _c_characterGenerator8x8[1078] = 8'h7e;
assign _c_characterGenerator8x8[1079] = 8'h00;
assign _c_characterGenerator8x8[1080] = 8'h00;
assign _c_characterGenerator8x8[1081] = 8'h00;
assign _c_characterGenerator8x8[1082] = 8'h78;
assign _c_characterGenerator8x8[1083] = 8'hc0;
assign _c_characterGenerator8x8[1084] = 8'hc0;
assign _c_characterGenerator8x8[1085] = 8'h78;
assign _c_characterGenerator8x8[1086] = 8'h0c;
assign _c_characterGenerator8x8[1087] = 8'h38;
assign _c_characterGenerator8x8[1088] = 8'h7e;
assign _c_characterGenerator8x8[1089] = 8'hc3;
assign _c_characterGenerator8x8[1090] = 8'h3c;
assign _c_characterGenerator8x8[1091] = 8'h66;
assign _c_characterGenerator8x8[1092] = 8'h7e;
assign _c_characterGenerator8x8[1093] = 8'h60;
assign _c_characterGenerator8x8[1094] = 8'h3c;
assign _c_characterGenerator8x8[1095] = 8'h00;
assign _c_characterGenerator8x8[1096] = 8'hcc;
assign _c_characterGenerator8x8[1097] = 8'h00;
assign _c_characterGenerator8x8[1098] = 8'h78;
assign _c_characterGenerator8x8[1099] = 8'hcc;
assign _c_characterGenerator8x8[1100] = 8'hfc;
assign _c_characterGenerator8x8[1101] = 8'hc0;
assign _c_characterGenerator8x8[1102] = 8'h78;
assign _c_characterGenerator8x8[1103] = 8'h00;
assign _c_characterGenerator8x8[1104] = 8'he0;
assign _c_characterGenerator8x8[1105] = 8'h00;
assign _c_characterGenerator8x8[1106] = 8'h78;
assign _c_characterGenerator8x8[1107] = 8'hcc;
assign _c_characterGenerator8x8[1108] = 8'hfc;
assign _c_characterGenerator8x8[1109] = 8'hc0;
assign _c_characterGenerator8x8[1110] = 8'h78;
assign _c_characterGenerator8x8[1111] = 8'h00;
assign _c_characterGenerator8x8[1112] = 8'hcc;
assign _c_characterGenerator8x8[1113] = 8'h00;
assign _c_characterGenerator8x8[1114] = 8'h70;
assign _c_characterGenerator8x8[1115] = 8'h30;
assign _c_characterGenerator8x8[1116] = 8'h30;
assign _c_characterGenerator8x8[1117] = 8'h30;
assign _c_characterGenerator8x8[1118] = 8'h78;
assign _c_characterGenerator8x8[1119] = 8'h00;
assign _c_characterGenerator8x8[1120] = 8'h7c;
assign _c_characterGenerator8x8[1121] = 8'hc6;
assign _c_characterGenerator8x8[1122] = 8'h38;
assign _c_characterGenerator8x8[1123] = 8'h18;
assign _c_characterGenerator8x8[1124] = 8'h18;
assign _c_characterGenerator8x8[1125] = 8'h18;
assign _c_characterGenerator8x8[1126] = 8'h3c;
assign _c_characterGenerator8x8[1127] = 8'h00;
assign _c_characterGenerator8x8[1128] = 8'he0;
assign _c_characterGenerator8x8[1129] = 8'h00;
assign _c_characterGenerator8x8[1130] = 8'h70;
assign _c_characterGenerator8x8[1131] = 8'h30;
assign _c_characterGenerator8x8[1132] = 8'h30;
assign _c_characterGenerator8x8[1133] = 8'h30;
assign _c_characterGenerator8x8[1134] = 8'h78;
assign _c_characterGenerator8x8[1135] = 8'h00;
assign _c_characterGenerator8x8[1136] = 8'hc6;
assign _c_characterGenerator8x8[1137] = 8'h38;
assign _c_characterGenerator8x8[1138] = 8'h6c;
assign _c_characterGenerator8x8[1139] = 8'hc6;
assign _c_characterGenerator8x8[1140] = 8'hfe;
assign _c_characterGenerator8x8[1141] = 8'hc6;
assign _c_characterGenerator8x8[1142] = 8'hc6;
assign _c_characterGenerator8x8[1143] = 8'h00;
assign _c_characterGenerator8x8[1144] = 8'h30;
assign _c_characterGenerator8x8[1145] = 8'h30;
assign _c_characterGenerator8x8[1146] = 8'h00;
assign _c_characterGenerator8x8[1147] = 8'h78;
assign _c_characterGenerator8x8[1148] = 8'hcc;
assign _c_characterGenerator8x8[1149] = 8'hfc;
assign _c_characterGenerator8x8[1150] = 8'hcc;
assign _c_characterGenerator8x8[1151] = 8'h00;
assign _c_characterGenerator8x8[1152] = 8'h1c;
assign _c_characterGenerator8x8[1153] = 8'h00;
assign _c_characterGenerator8x8[1154] = 8'hfc;
assign _c_characterGenerator8x8[1155] = 8'h60;
assign _c_characterGenerator8x8[1156] = 8'h78;
assign _c_characterGenerator8x8[1157] = 8'h60;
assign _c_characterGenerator8x8[1158] = 8'hfc;
assign _c_characterGenerator8x8[1159] = 8'h00;
assign _c_characterGenerator8x8[1160] = 8'h00;
assign _c_characterGenerator8x8[1161] = 8'h00;
assign _c_characterGenerator8x8[1162] = 8'h7f;
assign _c_characterGenerator8x8[1163] = 8'h0c;
assign _c_characterGenerator8x8[1164] = 8'h7f;
assign _c_characterGenerator8x8[1165] = 8'hcc;
assign _c_characterGenerator8x8[1166] = 8'h7f;
assign _c_characterGenerator8x8[1167] = 8'h00;
assign _c_characterGenerator8x8[1168] = 8'h3e;
assign _c_characterGenerator8x8[1169] = 8'h6c;
assign _c_characterGenerator8x8[1170] = 8'hcc;
assign _c_characterGenerator8x8[1171] = 8'hfe;
assign _c_characterGenerator8x8[1172] = 8'hcc;
assign _c_characterGenerator8x8[1173] = 8'hcc;
assign _c_characterGenerator8x8[1174] = 8'hce;
assign _c_characterGenerator8x8[1175] = 8'h00;
assign _c_characterGenerator8x8[1176] = 8'h78;
assign _c_characterGenerator8x8[1177] = 8'hcc;
assign _c_characterGenerator8x8[1178] = 8'h00;
assign _c_characterGenerator8x8[1179] = 8'h78;
assign _c_characterGenerator8x8[1180] = 8'hcc;
assign _c_characterGenerator8x8[1181] = 8'hcc;
assign _c_characterGenerator8x8[1182] = 8'h78;
assign _c_characterGenerator8x8[1183] = 8'h00;
assign _c_characterGenerator8x8[1184] = 8'h00;
assign _c_characterGenerator8x8[1185] = 8'hcc;
assign _c_characterGenerator8x8[1186] = 8'h00;
assign _c_characterGenerator8x8[1187] = 8'h78;
assign _c_characterGenerator8x8[1188] = 8'hcc;
assign _c_characterGenerator8x8[1189] = 8'hcc;
assign _c_characterGenerator8x8[1190] = 8'h78;
assign _c_characterGenerator8x8[1191] = 8'h00;
assign _c_characterGenerator8x8[1192] = 8'h00;
assign _c_characterGenerator8x8[1193] = 8'he0;
assign _c_characterGenerator8x8[1194] = 8'h00;
assign _c_characterGenerator8x8[1195] = 8'h78;
assign _c_characterGenerator8x8[1196] = 8'hcc;
assign _c_characterGenerator8x8[1197] = 8'hcc;
assign _c_characterGenerator8x8[1198] = 8'h78;
assign _c_characterGenerator8x8[1199] = 8'h00;
assign _c_characterGenerator8x8[1200] = 8'h78;
assign _c_characterGenerator8x8[1201] = 8'hcc;
assign _c_characterGenerator8x8[1202] = 8'h00;
assign _c_characterGenerator8x8[1203] = 8'hcc;
assign _c_characterGenerator8x8[1204] = 8'hcc;
assign _c_characterGenerator8x8[1205] = 8'hcc;
assign _c_characterGenerator8x8[1206] = 8'h7e;
assign _c_characterGenerator8x8[1207] = 8'h00;
assign _c_characterGenerator8x8[1208] = 8'h00;
assign _c_characterGenerator8x8[1209] = 8'he0;
assign _c_characterGenerator8x8[1210] = 8'h00;
assign _c_characterGenerator8x8[1211] = 8'hcc;
assign _c_characterGenerator8x8[1212] = 8'hcc;
assign _c_characterGenerator8x8[1213] = 8'hcc;
assign _c_characterGenerator8x8[1214] = 8'h7e;
assign _c_characterGenerator8x8[1215] = 8'h00;
assign _c_characterGenerator8x8[1216] = 8'h00;
assign _c_characterGenerator8x8[1217] = 8'hcc;
assign _c_characterGenerator8x8[1218] = 8'h00;
assign _c_characterGenerator8x8[1219] = 8'hcc;
assign _c_characterGenerator8x8[1220] = 8'hcc;
assign _c_characterGenerator8x8[1221] = 8'h7c;
assign _c_characterGenerator8x8[1222] = 8'h0c;
assign _c_characterGenerator8x8[1223] = 8'hf8;
assign _c_characterGenerator8x8[1224] = 8'hc3;
assign _c_characterGenerator8x8[1225] = 8'h18;
assign _c_characterGenerator8x8[1226] = 8'h3c;
assign _c_characterGenerator8x8[1227] = 8'h66;
assign _c_characterGenerator8x8[1228] = 8'h66;
assign _c_characterGenerator8x8[1229] = 8'h3c;
assign _c_characterGenerator8x8[1230] = 8'h18;
assign _c_characterGenerator8x8[1231] = 8'h00;
assign _c_characterGenerator8x8[1232] = 8'hcc;
assign _c_characterGenerator8x8[1233] = 8'h00;
assign _c_characterGenerator8x8[1234] = 8'hcc;
assign _c_characterGenerator8x8[1235] = 8'hcc;
assign _c_characterGenerator8x8[1236] = 8'hcc;
assign _c_characterGenerator8x8[1237] = 8'hcc;
assign _c_characterGenerator8x8[1238] = 8'h78;
assign _c_characterGenerator8x8[1239] = 8'h00;
assign _c_characterGenerator8x8[1240] = 8'h18;
assign _c_characterGenerator8x8[1241] = 8'h18;
assign _c_characterGenerator8x8[1242] = 8'h7e;
assign _c_characterGenerator8x8[1243] = 8'hc0;
assign _c_characterGenerator8x8[1244] = 8'hc0;
assign _c_characterGenerator8x8[1245] = 8'h7e;
assign _c_characterGenerator8x8[1246] = 8'h18;
assign _c_characterGenerator8x8[1247] = 8'h18;
assign _c_characterGenerator8x8[1248] = 8'h38;
assign _c_characterGenerator8x8[1249] = 8'h6c;
assign _c_characterGenerator8x8[1250] = 8'h64;
assign _c_characterGenerator8x8[1251] = 8'hf0;
assign _c_characterGenerator8x8[1252] = 8'h60;
assign _c_characterGenerator8x8[1253] = 8'he6;
assign _c_characterGenerator8x8[1254] = 8'hfc;
assign _c_characterGenerator8x8[1255] = 8'h00;
assign _c_characterGenerator8x8[1256] = 8'hcc;
assign _c_characterGenerator8x8[1257] = 8'hcc;
assign _c_characterGenerator8x8[1258] = 8'h78;
assign _c_characterGenerator8x8[1259] = 8'hfc;
assign _c_characterGenerator8x8[1260] = 8'h30;
assign _c_characterGenerator8x8[1261] = 8'hfc;
assign _c_characterGenerator8x8[1262] = 8'h30;
assign _c_characterGenerator8x8[1263] = 8'h30;
assign _c_characterGenerator8x8[1264] = 8'hf8;
assign _c_characterGenerator8x8[1265] = 8'hcc;
assign _c_characterGenerator8x8[1266] = 8'hcc;
assign _c_characterGenerator8x8[1267] = 8'hfa;
assign _c_characterGenerator8x8[1268] = 8'hc6;
assign _c_characterGenerator8x8[1269] = 8'hcf;
assign _c_characterGenerator8x8[1270] = 8'hc6;
assign _c_characterGenerator8x8[1271] = 8'hc7;
assign _c_characterGenerator8x8[1272] = 8'h0e;
assign _c_characterGenerator8x8[1273] = 8'h1b;
assign _c_characterGenerator8x8[1274] = 8'h18;
assign _c_characterGenerator8x8[1275] = 8'h3c;
assign _c_characterGenerator8x8[1276] = 8'h18;
assign _c_characterGenerator8x8[1277] = 8'h18;
assign _c_characterGenerator8x8[1278] = 8'hd8;
assign _c_characterGenerator8x8[1279] = 8'h70;
assign _c_characterGenerator8x8[1280] = 8'h1c;
assign _c_characterGenerator8x8[1281] = 8'h00;
assign _c_characterGenerator8x8[1282] = 8'h78;
assign _c_characterGenerator8x8[1283] = 8'h0c;
assign _c_characterGenerator8x8[1284] = 8'h7c;
assign _c_characterGenerator8x8[1285] = 8'hcc;
assign _c_characterGenerator8x8[1286] = 8'h7e;
assign _c_characterGenerator8x8[1287] = 8'h00;
assign _c_characterGenerator8x8[1288] = 8'h38;
assign _c_characterGenerator8x8[1289] = 8'h00;
assign _c_characterGenerator8x8[1290] = 8'h70;
assign _c_characterGenerator8x8[1291] = 8'h30;
assign _c_characterGenerator8x8[1292] = 8'h30;
assign _c_characterGenerator8x8[1293] = 8'h30;
assign _c_characterGenerator8x8[1294] = 8'h78;
assign _c_characterGenerator8x8[1295] = 8'h00;
assign _c_characterGenerator8x8[1296] = 8'h00;
assign _c_characterGenerator8x8[1297] = 8'h1c;
assign _c_characterGenerator8x8[1298] = 8'h00;
assign _c_characterGenerator8x8[1299] = 8'h78;
assign _c_characterGenerator8x8[1300] = 8'hcc;
assign _c_characterGenerator8x8[1301] = 8'hcc;
assign _c_characterGenerator8x8[1302] = 8'h78;
assign _c_characterGenerator8x8[1303] = 8'h00;
assign _c_characterGenerator8x8[1304] = 8'h00;
assign _c_characterGenerator8x8[1305] = 8'h1c;
assign _c_characterGenerator8x8[1306] = 8'h00;
assign _c_characterGenerator8x8[1307] = 8'hcc;
assign _c_characterGenerator8x8[1308] = 8'hcc;
assign _c_characterGenerator8x8[1309] = 8'hcc;
assign _c_characterGenerator8x8[1310] = 8'h7e;
assign _c_characterGenerator8x8[1311] = 8'h00;
assign _c_characterGenerator8x8[1312] = 8'h00;
assign _c_characterGenerator8x8[1313] = 8'hf8;
assign _c_characterGenerator8x8[1314] = 8'h00;
assign _c_characterGenerator8x8[1315] = 8'hf8;
assign _c_characterGenerator8x8[1316] = 8'hcc;
assign _c_characterGenerator8x8[1317] = 8'hcc;
assign _c_characterGenerator8x8[1318] = 8'hcc;
assign _c_characterGenerator8x8[1319] = 8'h00;
assign _c_characterGenerator8x8[1320] = 8'hfc;
assign _c_characterGenerator8x8[1321] = 8'h00;
assign _c_characterGenerator8x8[1322] = 8'hcc;
assign _c_characterGenerator8x8[1323] = 8'hec;
assign _c_characterGenerator8x8[1324] = 8'hfc;
assign _c_characterGenerator8x8[1325] = 8'hdc;
assign _c_characterGenerator8x8[1326] = 8'hcc;
assign _c_characterGenerator8x8[1327] = 8'h00;
assign _c_characterGenerator8x8[1328] = 8'h3c;
assign _c_characterGenerator8x8[1329] = 8'h6c;
assign _c_characterGenerator8x8[1330] = 8'h6c;
assign _c_characterGenerator8x8[1331] = 8'h3e;
assign _c_characterGenerator8x8[1332] = 8'h00;
assign _c_characterGenerator8x8[1333] = 8'h7e;
assign _c_characterGenerator8x8[1334] = 8'h00;
assign _c_characterGenerator8x8[1335] = 8'h00;
assign _c_characterGenerator8x8[1336] = 8'h38;
assign _c_characterGenerator8x8[1337] = 8'h6c;
assign _c_characterGenerator8x8[1338] = 8'h6c;
assign _c_characterGenerator8x8[1339] = 8'h38;
assign _c_characterGenerator8x8[1340] = 8'h00;
assign _c_characterGenerator8x8[1341] = 8'h7c;
assign _c_characterGenerator8x8[1342] = 8'h00;
assign _c_characterGenerator8x8[1343] = 8'h00;
assign _c_characterGenerator8x8[1344] = 8'h30;
assign _c_characterGenerator8x8[1345] = 8'h00;
assign _c_characterGenerator8x8[1346] = 8'h30;
assign _c_characterGenerator8x8[1347] = 8'h60;
assign _c_characterGenerator8x8[1348] = 8'hc0;
assign _c_characterGenerator8x8[1349] = 8'hcc;
assign _c_characterGenerator8x8[1350] = 8'h78;
assign _c_characterGenerator8x8[1351] = 8'h00;
assign _c_characterGenerator8x8[1352] = 8'h00;
assign _c_characterGenerator8x8[1353] = 8'h00;
assign _c_characterGenerator8x8[1354] = 8'h00;
assign _c_characterGenerator8x8[1355] = 8'hfc;
assign _c_characterGenerator8x8[1356] = 8'hc0;
assign _c_characterGenerator8x8[1357] = 8'hc0;
assign _c_characterGenerator8x8[1358] = 8'h00;
assign _c_characterGenerator8x8[1359] = 8'h00;
assign _c_characterGenerator8x8[1360] = 8'h00;
assign _c_characterGenerator8x8[1361] = 8'h00;
assign _c_characterGenerator8x8[1362] = 8'h00;
assign _c_characterGenerator8x8[1363] = 8'hfc;
assign _c_characterGenerator8x8[1364] = 8'h0c;
assign _c_characterGenerator8x8[1365] = 8'h0c;
assign _c_characterGenerator8x8[1366] = 8'h00;
assign _c_characterGenerator8x8[1367] = 8'h00;
assign _c_characterGenerator8x8[1368] = 8'hc3;
assign _c_characterGenerator8x8[1369] = 8'hc6;
assign _c_characterGenerator8x8[1370] = 8'hcc;
assign _c_characterGenerator8x8[1371] = 8'hde;
assign _c_characterGenerator8x8[1372] = 8'h33;
assign _c_characterGenerator8x8[1373] = 8'h66;
assign _c_characterGenerator8x8[1374] = 8'hcc;
assign _c_characterGenerator8x8[1375] = 8'h0f;
assign _c_characterGenerator8x8[1376] = 8'hc3;
assign _c_characterGenerator8x8[1377] = 8'hc6;
assign _c_characterGenerator8x8[1378] = 8'hcc;
assign _c_characterGenerator8x8[1379] = 8'hdb;
assign _c_characterGenerator8x8[1380] = 8'h37;
assign _c_characterGenerator8x8[1381] = 8'h6f;
assign _c_characterGenerator8x8[1382] = 8'hcf;
assign _c_characterGenerator8x8[1383] = 8'h03;
assign _c_characterGenerator8x8[1384] = 8'h18;
assign _c_characterGenerator8x8[1385] = 8'h18;
assign _c_characterGenerator8x8[1386] = 8'h00;
assign _c_characterGenerator8x8[1387] = 8'h18;
assign _c_characterGenerator8x8[1388] = 8'h18;
assign _c_characterGenerator8x8[1389] = 8'h18;
assign _c_characterGenerator8x8[1390] = 8'h18;
assign _c_characterGenerator8x8[1391] = 8'h00;
assign _c_characterGenerator8x8[1392] = 8'h00;
assign _c_characterGenerator8x8[1393] = 8'h33;
assign _c_characterGenerator8x8[1394] = 8'h66;
assign _c_characterGenerator8x8[1395] = 8'hcc;
assign _c_characterGenerator8x8[1396] = 8'h66;
assign _c_characterGenerator8x8[1397] = 8'h33;
assign _c_characterGenerator8x8[1398] = 8'h00;
assign _c_characterGenerator8x8[1399] = 8'h00;
assign _c_characterGenerator8x8[1400] = 8'h00;
assign _c_characterGenerator8x8[1401] = 8'hcc;
assign _c_characterGenerator8x8[1402] = 8'h66;
assign _c_characterGenerator8x8[1403] = 8'h33;
assign _c_characterGenerator8x8[1404] = 8'h66;
assign _c_characterGenerator8x8[1405] = 8'hcc;
assign _c_characterGenerator8x8[1406] = 8'h00;
assign _c_characterGenerator8x8[1407] = 8'h00;
assign _c_characterGenerator8x8[1408] = 8'h22;
assign _c_characterGenerator8x8[1409] = 8'h88;
assign _c_characterGenerator8x8[1410] = 8'h22;
assign _c_characterGenerator8x8[1411] = 8'h88;
assign _c_characterGenerator8x8[1412] = 8'h22;
assign _c_characterGenerator8x8[1413] = 8'h88;
assign _c_characterGenerator8x8[1414] = 8'h22;
assign _c_characterGenerator8x8[1415] = 8'h88;
assign _c_characterGenerator8x8[1416] = 8'h55;
assign _c_characterGenerator8x8[1417] = 8'haa;
assign _c_characterGenerator8x8[1418] = 8'h55;
assign _c_characterGenerator8x8[1419] = 8'haa;
assign _c_characterGenerator8x8[1420] = 8'h55;
assign _c_characterGenerator8x8[1421] = 8'haa;
assign _c_characterGenerator8x8[1422] = 8'h55;
assign _c_characterGenerator8x8[1423] = 8'haa;
assign _c_characterGenerator8x8[1424] = 8'hdb;
assign _c_characterGenerator8x8[1425] = 8'h77;
assign _c_characterGenerator8x8[1426] = 8'hdb;
assign _c_characterGenerator8x8[1427] = 8'hee;
assign _c_characterGenerator8x8[1428] = 8'hdb;
assign _c_characterGenerator8x8[1429] = 8'h77;
assign _c_characterGenerator8x8[1430] = 8'hdb;
assign _c_characterGenerator8x8[1431] = 8'hee;
assign _c_characterGenerator8x8[1432] = 8'h18;
assign _c_characterGenerator8x8[1433] = 8'h18;
assign _c_characterGenerator8x8[1434] = 8'h18;
assign _c_characterGenerator8x8[1435] = 8'h18;
assign _c_characterGenerator8x8[1436] = 8'h18;
assign _c_characterGenerator8x8[1437] = 8'h18;
assign _c_characterGenerator8x8[1438] = 8'h18;
assign _c_characterGenerator8x8[1439] = 8'h18;
assign _c_characterGenerator8x8[1440] = 8'h18;
assign _c_characterGenerator8x8[1441] = 8'h18;
assign _c_characterGenerator8x8[1442] = 8'h18;
assign _c_characterGenerator8x8[1443] = 8'h18;
assign _c_characterGenerator8x8[1444] = 8'hf8;
assign _c_characterGenerator8x8[1445] = 8'h18;
assign _c_characterGenerator8x8[1446] = 8'h18;
assign _c_characterGenerator8x8[1447] = 8'h18;
assign _c_characterGenerator8x8[1448] = 8'h18;
assign _c_characterGenerator8x8[1449] = 8'h18;
assign _c_characterGenerator8x8[1450] = 8'hf8;
assign _c_characterGenerator8x8[1451] = 8'h18;
assign _c_characterGenerator8x8[1452] = 8'hf8;
assign _c_characterGenerator8x8[1453] = 8'h18;
assign _c_characterGenerator8x8[1454] = 8'h18;
assign _c_characterGenerator8x8[1455] = 8'h18;
assign _c_characterGenerator8x8[1456] = 8'h36;
assign _c_characterGenerator8x8[1457] = 8'h36;
assign _c_characterGenerator8x8[1458] = 8'h36;
assign _c_characterGenerator8x8[1459] = 8'h36;
assign _c_characterGenerator8x8[1460] = 8'hf6;
assign _c_characterGenerator8x8[1461] = 8'h36;
assign _c_characterGenerator8x8[1462] = 8'h36;
assign _c_characterGenerator8x8[1463] = 8'h36;
assign _c_characterGenerator8x8[1464] = 8'h00;
assign _c_characterGenerator8x8[1465] = 8'h00;
assign _c_characterGenerator8x8[1466] = 8'h00;
assign _c_characterGenerator8x8[1467] = 8'h00;
assign _c_characterGenerator8x8[1468] = 8'hfe;
assign _c_characterGenerator8x8[1469] = 8'h36;
assign _c_characterGenerator8x8[1470] = 8'h36;
assign _c_characterGenerator8x8[1471] = 8'h36;
assign _c_characterGenerator8x8[1472] = 8'h00;
assign _c_characterGenerator8x8[1473] = 8'h00;
assign _c_characterGenerator8x8[1474] = 8'hf8;
assign _c_characterGenerator8x8[1475] = 8'h18;
assign _c_characterGenerator8x8[1476] = 8'hf8;
assign _c_characterGenerator8x8[1477] = 8'h18;
assign _c_characterGenerator8x8[1478] = 8'h18;
assign _c_characterGenerator8x8[1479] = 8'h18;
assign _c_characterGenerator8x8[1480] = 8'h36;
assign _c_characterGenerator8x8[1481] = 8'h36;
assign _c_characterGenerator8x8[1482] = 8'hf6;
assign _c_characterGenerator8x8[1483] = 8'h06;
assign _c_characterGenerator8x8[1484] = 8'hf6;
assign _c_characterGenerator8x8[1485] = 8'h36;
assign _c_characterGenerator8x8[1486] = 8'h36;
assign _c_characterGenerator8x8[1487] = 8'h36;
assign _c_characterGenerator8x8[1488] = 8'h36;
assign _c_characterGenerator8x8[1489] = 8'h36;
assign _c_characterGenerator8x8[1490] = 8'h36;
assign _c_characterGenerator8x8[1491] = 8'h36;
assign _c_characterGenerator8x8[1492] = 8'h36;
assign _c_characterGenerator8x8[1493] = 8'h36;
assign _c_characterGenerator8x8[1494] = 8'h36;
assign _c_characterGenerator8x8[1495] = 8'h36;
assign _c_characterGenerator8x8[1496] = 8'h00;
assign _c_characterGenerator8x8[1497] = 8'h00;
assign _c_characterGenerator8x8[1498] = 8'hfe;
assign _c_characterGenerator8x8[1499] = 8'h06;
assign _c_characterGenerator8x8[1500] = 8'hf6;
assign _c_characterGenerator8x8[1501] = 8'h36;
assign _c_characterGenerator8x8[1502] = 8'h36;
assign _c_characterGenerator8x8[1503] = 8'h36;
assign _c_characterGenerator8x8[1504] = 8'h36;
assign _c_characterGenerator8x8[1505] = 8'h36;
assign _c_characterGenerator8x8[1506] = 8'hf6;
assign _c_characterGenerator8x8[1507] = 8'h06;
assign _c_characterGenerator8x8[1508] = 8'hfe;
assign _c_characterGenerator8x8[1509] = 8'h00;
assign _c_characterGenerator8x8[1510] = 8'h00;
assign _c_characterGenerator8x8[1511] = 8'h00;
assign _c_characterGenerator8x8[1512] = 8'h36;
assign _c_characterGenerator8x8[1513] = 8'h36;
assign _c_characterGenerator8x8[1514] = 8'h36;
assign _c_characterGenerator8x8[1515] = 8'h36;
assign _c_characterGenerator8x8[1516] = 8'hfe;
assign _c_characterGenerator8x8[1517] = 8'h00;
assign _c_characterGenerator8x8[1518] = 8'h00;
assign _c_characterGenerator8x8[1519] = 8'h00;
assign _c_characterGenerator8x8[1520] = 8'h18;
assign _c_characterGenerator8x8[1521] = 8'h18;
assign _c_characterGenerator8x8[1522] = 8'hf8;
assign _c_characterGenerator8x8[1523] = 8'h18;
assign _c_characterGenerator8x8[1524] = 8'hf8;
assign _c_characterGenerator8x8[1525] = 8'h00;
assign _c_characterGenerator8x8[1526] = 8'h00;
assign _c_characterGenerator8x8[1527] = 8'h00;
assign _c_characterGenerator8x8[1528] = 8'h00;
assign _c_characterGenerator8x8[1529] = 8'h00;
assign _c_characterGenerator8x8[1530] = 8'h00;
assign _c_characterGenerator8x8[1531] = 8'h00;
assign _c_characterGenerator8x8[1532] = 8'hf8;
assign _c_characterGenerator8x8[1533] = 8'h18;
assign _c_characterGenerator8x8[1534] = 8'h18;
assign _c_characterGenerator8x8[1535] = 8'h18;
assign _c_characterGenerator8x8[1536] = 8'h18;
assign _c_characterGenerator8x8[1537] = 8'h18;
assign _c_characterGenerator8x8[1538] = 8'h18;
assign _c_characterGenerator8x8[1539] = 8'h18;
assign _c_characterGenerator8x8[1540] = 8'h1f;
assign _c_characterGenerator8x8[1541] = 8'h00;
assign _c_characterGenerator8x8[1542] = 8'h00;
assign _c_characterGenerator8x8[1543] = 8'h00;
assign _c_characterGenerator8x8[1544] = 8'h18;
assign _c_characterGenerator8x8[1545] = 8'h18;
assign _c_characterGenerator8x8[1546] = 8'h18;
assign _c_characterGenerator8x8[1547] = 8'h18;
assign _c_characterGenerator8x8[1548] = 8'hff;
assign _c_characterGenerator8x8[1549] = 8'h00;
assign _c_characterGenerator8x8[1550] = 8'h00;
assign _c_characterGenerator8x8[1551] = 8'h00;
assign _c_characterGenerator8x8[1552] = 8'h00;
assign _c_characterGenerator8x8[1553] = 8'h00;
assign _c_characterGenerator8x8[1554] = 8'h00;
assign _c_characterGenerator8x8[1555] = 8'h00;
assign _c_characterGenerator8x8[1556] = 8'hff;
assign _c_characterGenerator8x8[1557] = 8'h18;
assign _c_characterGenerator8x8[1558] = 8'h18;
assign _c_characterGenerator8x8[1559] = 8'h18;
assign _c_characterGenerator8x8[1560] = 8'h18;
assign _c_characterGenerator8x8[1561] = 8'h18;
assign _c_characterGenerator8x8[1562] = 8'h18;
assign _c_characterGenerator8x8[1563] = 8'h18;
assign _c_characterGenerator8x8[1564] = 8'h1f;
assign _c_characterGenerator8x8[1565] = 8'h18;
assign _c_characterGenerator8x8[1566] = 8'h18;
assign _c_characterGenerator8x8[1567] = 8'h18;
assign _c_characterGenerator8x8[1568] = 8'h00;
assign _c_characterGenerator8x8[1569] = 8'h00;
assign _c_characterGenerator8x8[1570] = 8'h00;
assign _c_characterGenerator8x8[1571] = 8'h00;
assign _c_characterGenerator8x8[1572] = 8'hff;
assign _c_characterGenerator8x8[1573] = 8'h00;
assign _c_characterGenerator8x8[1574] = 8'h00;
assign _c_characterGenerator8x8[1575] = 8'h00;
assign _c_characterGenerator8x8[1576] = 8'h18;
assign _c_characterGenerator8x8[1577] = 8'h18;
assign _c_characterGenerator8x8[1578] = 8'h18;
assign _c_characterGenerator8x8[1579] = 8'h18;
assign _c_characterGenerator8x8[1580] = 8'hff;
assign _c_characterGenerator8x8[1581] = 8'h18;
assign _c_characterGenerator8x8[1582] = 8'h18;
assign _c_characterGenerator8x8[1583] = 8'h18;
assign _c_characterGenerator8x8[1584] = 8'h18;
assign _c_characterGenerator8x8[1585] = 8'h18;
assign _c_characterGenerator8x8[1586] = 8'h1f;
assign _c_characterGenerator8x8[1587] = 8'h18;
assign _c_characterGenerator8x8[1588] = 8'h1f;
assign _c_characterGenerator8x8[1589] = 8'h18;
assign _c_characterGenerator8x8[1590] = 8'h18;
assign _c_characterGenerator8x8[1591] = 8'h18;
assign _c_characterGenerator8x8[1592] = 8'h36;
assign _c_characterGenerator8x8[1593] = 8'h36;
assign _c_characterGenerator8x8[1594] = 8'h36;
assign _c_characterGenerator8x8[1595] = 8'h36;
assign _c_characterGenerator8x8[1596] = 8'h37;
assign _c_characterGenerator8x8[1597] = 8'h36;
assign _c_characterGenerator8x8[1598] = 8'h36;
assign _c_characterGenerator8x8[1599] = 8'h36;
assign _c_characterGenerator8x8[1600] = 8'h36;
assign _c_characterGenerator8x8[1601] = 8'h36;
assign _c_characterGenerator8x8[1602] = 8'h37;
assign _c_characterGenerator8x8[1603] = 8'h30;
assign _c_characterGenerator8x8[1604] = 8'h3f;
assign _c_characterGenerator8x8[1605] = 8'h00;
assign _c_characterGenerator8x8[1606] = 8'h00;
assign _c_characterGenerator8x8[1607] = 8'h00;
assign _c_characterGenerator8x8[1608] = 8'h00;
assign _c_characterGenerator8x8[1609] = 8'h00;
assign _c_characterGenerator8x8[1610] = 8'h3f;
assign _c_characterGenerator8x8[1611] = 8'h30;
assign _c_characterGenerator8x8[1612] = 8'h37;
assign _c_characterGenerator8x8[1613] = 8'h36;
assign _c_characterGenerator8x8[1614] = 8'h36;
assign _c_characterGenerator8x8[1615] = 8'h36;
assign _c_characterGenerator8x8[1616] = 8'h36;
assign _c_characterGenerator8x8[1617] = 8'h36;
assign _c_characterGenerator8x8[1618] = 8'hf7;
assign _c_characterGenerator8x8[1619] = 8'h00;
assign _c_characterGenerator8x8[1620] = 8'hff;
assign _c_characterGenerator8x8[1621] = 8'h00;
assign _c_characterGenerator8x8[1622] = 8'h00;
assign _c_characterGenerator8x8[1623] = 8'h00;
assign _c_characterGenerator8x8[1624] = 8'h00;
assign _c_characterGenerator8x8[1625] = 8'h00;
assign _c_characterGenerator8x8[1626] = 8'hff;
assign _c_characterGenerator8x8[1627] = 8'h00;
assign _c_characterGenerator8x8[1628] = 8'hf7;
assign _c_characterGenerator8x8[1629] = 8'h36;
assign _c_characterGenerator8x8[1630] = 8'h36;
assign _c_characterGenerator8x8[1631] = 8'h36;
assign _c_characterGenerator8x8[1632] = 8'h36;
assign _c_characterGenerator8x8[1633] = 8'h36;
assign _c_characterGenerator8x8[1634] = 8'h37;
assign _c_characterGenerator8x8[1635] = 8'h30;
assign _c_characterGenerator8x8[1636] = 8'h37;
assign _c_characterGenerator8x8[1637] = 8'h36;
assign _c_characterGenerator8x8[1638] = 8'h36;
assign _c_characterGenerator8x8[1639] = 8'h36;
assign _c_characterGenerator8x8[1640] = 8'h00;
assign _c_characterGenerator8x8[1641] = 8'h00;
assign _c_characterGenerator8x8[1642] = 8'hff;
assign _c_characterGenerator8x8[1643] = 8'h00;
assign _c_characterGenerator8x8[1644] = 8'hff;
assign _c_characterGenerator8x8[1645] = 8'h00;
assign _c_characterGenerator8x8[1646] = 8'h00;
assign _c_characterGenerator8x8[1647] = 8'h00;
assign _c_characterGenerator8x8[1648] = 8'h36;
assign _c_characterGenerator8x8[1649] = 8'h36;
assign _c_characterGenerator8x8[1650] = 8'hf7;
assign _c_characterGenerator8x8[1651] = 8'h00;
assign _c_characterGenerator8x8[1652] = 8'hf7;
assign _c_characterGenerator8x8[1653] = 8'h36;
assign _c_characterGenerator8x8[1654] = 8'h36;
assign _c_characterGenerator8x8[1655] = 8'h36;
assign _c_characterGenerator8x8[1656] = 8'h18;
assign _c_characterGenerator8x8[1657] = 8'h18;
assign _c_characterGenerator8x8[1658] = 8'hff;
assign _c_characterGenerator8x8[1659] = 8'h00;
assign _c_characterGenerator8x8[1660] = 8'hff;
assign _c_characterGenerator8x8[1661] = 8'h00;
assign _c_characterGenerator8x8[1662] = 8'h00;
assign _c_characterGenerator8x8[1663] = 8'h00;
assign _c_characterGenerator8x8[1664] = 8'h36;
assign _c_characterGenerator8x8[1665] = 8'h36;
assign _c_characterGenerator8x8[1666] = 8'h36;
assign _c_characterGenerator8x8[1667] = 8'h36;
assign _c_characterGenerator8x8[1668] = 8'hff;
assign _c_characterGenerator8x8[1669] = 8'h00;
assign _c_characterGenerator8x8[1670] = 8'h00;
assign _c_characterGenerator8x8[1671] = 8'h00;
assign _c_characterGenerator8x8[1672] = 8'h00;
assign _c_characterGenerator8x8[1673] = 8'h00;
assign _c_characterGenerator8x8[1674] = 8'hff;
assign _c_characterGenerator8x8[1675] = 8'h00;
assign _c_characterGenerator8x8[1676] = 8'hff;
assign _c_characterGenerator8x8[1677] = 8'h18;
assign _c_characterGenerator8x8[1678] = 8'h18;
assign _c_characterGenerator8x8[1679] = 8'h18;
assign _c_characterGenerator8x8[1680] = 8'h00;
assign _c_characterGenerator8x8[1681] = 8'h00;
assign _c_characterGenerator8x8[1682] = 8'h00;
assign _c_characterGenerator8x8[1683] = 8'h00;
assign _c_characterGenerator8x8[1684] = 8'hff;
assign _c_characterGenerator8x8[1685] = 8'h36;
assign _c_characterGenerator8x8[1686] = 8'h36;
assign _c_characterGenerator8x8[1687] = 8'h36;
assign _c_characterGenerator8x8[1688] = 8'h36;
assign _c_characterGenerator8x8[1689] = 8'h36;
assign _c_characterGenerator8x8[1690] = 8'h36;
assign _c_characterGenerator8x8[1691] = 8'h36;
assign _c_characterGenerator8x8[1692] = 8'h3f;
assign _c_characterGenerator8x8[1693] = 8'h00;
assign _c_characterGenerator8x8[1694] = 8'h00;
assign _c_characterGenerator8x8[1695] = 8'h00;
assign _c_characterGenerator8x8[1696] = 8'h18;
assign _c_characterGenerator8x8[1697] = 8'h18;
assign _c_characterGenerator8x8[1698] = 8'h1f;
assign _c_characterGenerator8x8[1699] = 8'h18;
assign _c_characterGenerator8x8[1700] = 8'h1f;
assign _c_characterGenerator8x8[1701] = 8'h00;
assign _c_characterGenerator8x8[1702] = 8'h00;
assign _c_characterGenerator8x8[1703] = 8'h00;
assign _c_characterGenerator8x8[1704] = 8'h00;
assign _c_characterGenerator8x8[1705] = 8'h00;
assign _c_characterGenerator8x8[1706] = 8'h1f;
assign _c_characterGenerator8x8[1707] = 8'h18;
assign _c_characterGenerator8x8[1708] = 8'h1f;
assign _c_characterGenerator8x8[1709] = 8'h18;
assign _c_characterGenerator8x8[1710] = 8'h18;
assign _c_characterGenerator8x8[1711] = 8'h18;
assign _c_characterGenerator8x8[1712] = 8'h00;
assign _c_characterGenerator8x8[1713] = 8'h00;
assign _c_characterGenerator8x8[1714] = 8'h00;
assign _c_characterGenerator8x8[1715] = 8'h00;
assign _c_characterGenerator8x8[1716] = 8'h3f;
assign _c_characterGenerator8x8[1717] = 8'h36;
assign _c_characterGenerator8x8[1718] = 8'h36;
assign _c_characterGenerator8x8[1719] = 8'h36;
assign _c_characterGenerator8x8[1720] = 8'h36;
assign _c_characterGenerator8x8[1721] = 8'h36;
assign _c_characterGenerator8x8[1722] = 8'h36;
assign _c_characterGenerator8x8[1723] = 8'h36;
assign _c_characterGenerator8x8[1724] = 8'hff;
assign _c_characterGenerator8x8[1725] = 8'h36;
assign _c_characterGenerator8x8[1726] = 8'h36;
assign _c_characterGenerator8x8[1727] = 8'h36;
assign _c_characterGenerator8x8[1728] = 8'h18;
assign _c_characterGenerator8x8[1729] = 8'h18;
assign _c_characterGenerator8x8[1730] = 8'hff;
assign _c_characterGenerator8x8[1731] = 8'h18;
assign _c_characterGenerator8x8[1732] = 8'hff;
assign _c_characterGenerator8x8[1733] = 8'h18;
assign _c_characterGenerator8x8[1734] = 8'h18;
assign _c_characterGenerator8x8[1735] = 8'h18;
assign _c_characterGenerator8x8[1736] = 8'h18;
assign _c_characterGenerator8x8[1737] = 8'h18;
assign _c_characterGenerator8x8[1738] = 8'h18;
assign _c_characterGenerator8x8[1739] = 8'h18;
assign _c_characterGenerator8x8[1740] = 8'hf8;
assign _c_characterGenerator8x8[1741] = 8'h00;
assign _c_characterGenerator8x8[1742] = 8'h00;
assign _c_characterGenerator8x8[1743] = 8'h00;
assign _c_characterGenerator8x8[1744] = 8'h00;
assign _c_characterGenerator8x8[1745] = 8'h00;
assign _c_characterGenerator8x8[1746] = 8'h00;
assign _c_characterGenerator8x8[1747] = 8'h00;
assign _c_characterGenerator8x8[1748] = 8'h1f;
assign _c_characterGenerator8x8[1749] = 8'h18;
assign _c_characterGenerator8x8[1750] = 8'h18;
assign _c_characterGenerator8x8[1751] = 8'h18;
assign _c_characterGenerator8x8[1752] = 8'hff;
assign _c_characterGenerator8x8[1753] = 8'hff;
assign _c_characterGenerator8x8[1754] = 8'hff;
assign _c_characterGenerator8x8[1755] = 8'hff;
assign _c_characterGenerator8x8[1756] = 8'hff;
assign _c_characterGenerator8x8[1757] = 8'hff;
assign _c_characterGenerator8x8[1758] = 8'hff;
assign _c_characterGenerator8x8[1759] = 8'hff;
assign _c_characterGenerator8x8[1760] = 8'h00;
assign _c_characterGenerator8x8[1761] = 8'h00;
assign _c_characterGenerator8x8[1762] = 8'h00;
assign _c_characterGenerator8x8[1763] = 8'h00;
assign _c_characterGenerator8x8[1764] = 8'hff;
assign _c_characterGenerator8x8[1765] = 8'hff;
assign _c_characterGenerator8x8[1766] = 8'hff;
assign _c_characterGenerator8x8[1767] = 8'hff;
assign _c_characterGenerator8x8[1768] = 8'hf0;
assign _c_characterGenerator8x8[1769] = 8'hf0;
assign _c_characterGenerator8x8[1770] = 8'hf0;
assign _c_characterGenerator8x8[1771] = 8'hf0;
assign _c_characterGenerator8x8[1772] = 8'hf0;
assign _c_characterGenerator8x8[1773] = 8'hf0;
assign _c_characterGenerator8x8[1774] = 8'hf0;
assign _c_characterGenerator8x8[1775] = 8'hf0;
assign _c_characterGenerator8x8[1776] = 8'h0f;
assign _c_characterGenerator8x8[1777] = 8'h0f;
assign _c_characterGenerator8x8[1778] = 8'h0f;
assign _c_characterGenerator8x8[1779] = 8'h0f;
assign _c_characterGenerator8x8[1780] = 8'h0f;
assign _c_characterGenerator8x8[1781] = 8'h0f;
assign _c_characterGenerator8x8[1782] = 8'h0f;
assign _c_characterGenerator8x8[1783] = 8'h0f;
assign _c_characterGenerator8x8[1784] = 8'hff;
assign _c_characterGenerator8x8[1785] = 8'hff;
assign _c_characterGenerator8x8[1786] = 8'hff;
assign _c_characterGenerator8x8[1787] = 8'hff;
assign _c_characterGenerator8x8[1788] = 8'h00;
assign _c_characterGenerator8x8[1789] = 8'h00;
assign _c_characterGenerator8x8[1790] = 8'h00;
assign _c_characterGenerator8x8[1791] = 8'h00;
assign _c_characterGenerator8x8[1792] = 8'h00;
assign _c_characterGenerator8x8[1793] = 8'h00;
assign _c_characterGenerator8x8[1794] = 8'h76;
assign _c_characterGenerator8x8[1795] = 8'hdc;
assign _c_characterGenerator8x8[1796] = 8'hc8;
assign _c_characterGenerator8x8[1797] = 8'hdc;
assign _c_characterGenerator8x8[1798] = 8'h76;
assign _c_characterGenerator8x8[1799] = 8'h00;
assign _c_characterGenerator8x8[1800] = 8'h00;
assign _c_characterGenerator8x8[1801] = 8'h78;
assign _c_characterGenerator8x8[1802] = 8'hcc;
assign _c_characterGenerator8x8[1803] = 8'hf8;
assign _c_characterGenerator8x8[1804] = 8'hcc;
assign _c_characterGenerator8x8[1805] = 8'hf8;
assign _c_characterGenerator8x8[1806] = 8'hc0;
assign _c_characterGenerator8x8[1807] = 8'hc0;
assign _c_characterGenerator8x8[1808] = 8'h00;
assign _c_characterGenerator8x8[1809] = 8'hfc;
assign _c_characterGenerator8x8[1810] = 8'hcc;
assign _c_characterGenerator8x8[1811] = 8'hc0;
assign _c_characterGenerator8x8[1812] = 8'hc0;
assign _c_characterGenerator8x8[1813] = 8'hc0;
assign _c_characterGenerator8x8[1814] = 8'hc0;
assign _c_characterGenerator8x8[1815] = 8'h00;
assign _c_characterGenerator8x8[1816] = 8'h00;
assign _c_characterGenerator8x8[1817] = 8'hfe;
assign _c_characterGenerator8x8[1818] = 8'h6c;
assign _c_characterGenerator8x8[1819] = 8'h6c;
assign _c_characterGenerator8x8[1820] = 8'h6c;
assign _c_characterGenerator8x8[1821] = 8'h6c;
assign _c_characterGenerator8x8[1822] = 8'h6c;
assign _c_characterGenerator8x8[1823] = 8'h00;
assign _c_characterGenerator8x8[1824] = 8'hfc;
assign _c_characterGenerator8x8[1825] = 8'hcc;
assign _c_characterGenerator8x8[1826] = 8'h60;
assign _c_characterGenerator8x8[1827] = 8'h30;
assign _c_characterGenerator8x8[1828] = 8'h60;
assign _c_characterGenerator8x8[1829] = 8'hcc;
assign _c_characterGenerator8x8[1830] = 8'hfc;
assign _c_characterGenerator8x8[1831] = 8'h00;
assign _c_characterGenerator8x8[1832] = 8'h00;
assign _c_characterGenerator8x8[1833] = 8'h00;
assign _c_characterGenerator8x8[1834] = 8'h7e;
assign _c_characterGenerator8x8[1835] = 8'hd8;
assign _c_characterGenerator8x8[1836] = 8'hd8;
assign _c_characterGenerator8x8[1837] = 8'hd8;
assign _c_characterGenerator8x8[1838] = 8'h70;
assign _c_characterGenerator8x8[1839] = 8'h00;
assign _c_characterGenerator8x8[1840] = 8'h00;
assign _c_characterGenerator8x8[1841] = 8'h66;
assign _c_characterGenerator8x8[1842] = 8'h66;
assign _c_characterGenerator8x8[1843] = 8'h66;
assign _c_characterGenerator8x8[1844] = 8'h66;
assign _c_characterGenerator8x8[1845] = 8'h7c;
assign _c_characterGenerator8x8[1846] = 8'h60;
assign _c_characterGenerator8x8[1847] = 8'hc0;
assign _c_characterGenerator8x8[1848] = 8'h00;
assign _c_characterGenerator8x8[1849] = 8'h76;
assign _c_characterGenerator8x8[1850] = 8'hdc;
assign _c_characterGenerator8x8[1851] = 8'h18;
assign _c_characterGenerator8x8[1852] = 8'h18;
assign _c_characterGenerator8x8[1853] = 8'h18;
assign _c_characterGenerator8x8[1854] = 8'h18;
assign _c_characterGenerator8x8[1855] = 8'h00;
assign _c_characterGenerator8x8[1856] = 8'hfc;
assign _c_characterGenerator8x8[1857] = 8'h30;
assign _c_characterGenerator8x8[1858] = 8'h78;
assign _c_characterGenerator8x8[1859] = 8'hcc;
assign _c_characterGenerator8x8[1860] = 8'hcc;
assign _c_characterGenerator8x8[1861] = 8'h78;
assign _c_characterGenerator8x8[1862] = 8'h30;
assign _c_characterGenerator8x8[1863] = 8'hfc;
assign _c_characterGenerator8x8[1864] = 8'h38;
assign _c_characterGenerator8x8[1865] = 8'h6c;
assign _c_characterGenerator8x8[1866] = 8'hc6;
assign _c_characterGenerator8x8[1867] = 8'hfe;
assign _c_characterGenerator8x8[1868] = 8'hc6;
assign _c_characterGenerator8x8[1869] = 8'h6c;
assign _c_characterGenerator8x8[1870] = 8'h38;
assign _c_characterGenerator8x8[1871] = 8'h00;
assign _c_characterGenerator8x8[1872] = 8'h38;
assign _c_characterGenerator8x8[1873] = 8'h6c;
assign _c_characterGenerator8x8[1874] = 8'hc6;
assign _c_characterGenerator8x8[1875] = 8'hc6;
assign _c_characterGenerator8x8[1876] = 8'h6c;
assign _c_characterGenerator8x8[1877] = 8'h6c;
assign _c_characterGenerator8x8[1878] = 8'hee;
assign _c_characterGenerator8x8[1879] = 8'h00;
assign _c_characterGenerator8x8[1880] = 8'h1c;
assign _c_characterGenerator8x8[1881] = 8'h30;
assign _c_characterGenerator8x8[1882] = 8'h18;
assign _c_characterGenerator8x8[1883] = 8'h7c;
assign _c_characterGenerator8x8[1884] = 8'hcc;
assign _c_characterGenerator8x8[1885] = 8'hcc;
assign _c_characterGenerator8x8[1886] = 8'h78;
assign _c_characterGenerator8x8[1887] = 8'h00;
assign _c_characterGenerator8x8[1888] = 8'h00;
assign _c_characterGenerator8x8[1889] = 8'h00;
assign _c_characterGenerator8x8[1890] = 8'h7e;
assign _c_characterGenerator8x8[1891] = 8'hdb;
assign _c_characterGenerator8x8[1892] = 8'hdb;
assign _c_characterGenerator8x8[1893] = 8'h7e;
assign _c_characterGenerator8x8[1894] = 8'h00;
assign _c_characterGenerator8x8[1895] = 8'h00;
assign _c_characterGenerator8x8[1896] = 8'h06;
assign _c_characterGenerator8x8[1897] = 8'h0c;
assign _c_characterGenerator8x8[1898] = 8'h7e;
assign _c_characterGenerator8x8[1899] = 8'hdb;
assign _c_characterGenerator8x8[1900] = 8'hdb;
assign _c_characterGenerator8x8[1901] = 8'h7e;
assign _c_characterGenerator8x8[1902] = 8'h60;
assign _c_characterGenerator8x8[1903] = 8'hc0;
assign _c_characterGenerator8x8[1904] = 8'h38;
assign _c_characterGenerator8x8[1905] = 8'h60;
assign _c_characterGenerator8x8[1906] = 8'hc0;
assign _c_characterGenerator8x8[1907] = 8'hf8;
assign _c_characterGenerator8x8[1908] = 8'hc0;
assign _c_characterGenerator8x8[1909] = 8'h60;
assign _c_characterGenerator8x8[1910] = 8'h38;
assign _c_characterGenerator8x8[1911] = 8'h00;
assign _c_characterGenerator8x8[1912] = 8'h78;
assign _c_characterGenerator8x8[1913] = 8'hcc;
assign _c_characterGenerator8x8[1914] = 8'hcc;
assign _c_characterGenerator8x8[1915] = 8'hcc;
assign _c_characterGenerator8x8[1916] = 8'hcc;
assign _c_characterGenerator8x8[1917] = 8'hcc;
assign _c_characterGenerator8x8[1918] = 8'hcc;
assign _c_characterGenerator8x8[1919] = 8'h00;
assign _c_characterGenerator8x8[1920] = 8'h00;
assign _c_characterGenerator8x8[1921] = 8'hfc;
assign _c_characterGenerator8x8[1922] = 8'h00;
assign _c_characterGenerator8x8[1923] = 8'hfc;
assign _c_characterGenerator8x8[1924] = 8'h00;
assign _c_characterGenerator8x8[1925] = 8'hfc;
assign _c_characterGenerator8x8[1926] = 8'h00;
assign _c_characterGenerator8x8[1927] = 8'h00;
assign _c_characterGenerator8x8[1928] = 8'h30;
assign _c_characterGenerator8x8[1929] = 8'h30;
assign _c_characterGenerator8x8[1930] = 8'hfc;
assign _c_characterGenerator8x8[1931] = 8'h30;
assign _c_characterGenerator8x8[1932] = 8'h30;
assign _c_characterGenerator8x8[1933] = 8'h00;
assign _c_characterGenerator8x8[1934] = 8'hfc;
assign _c_characterGenerator8x8[1935] = 8'h00;
assign _c_characterGenerator8x8[1936] = 8'h60;
assign _c_characterGenerator8x8[1937] = 8'h30;
assign _c_characterGenerator8x8[1938] = 8'h18;
assign _c_characterGenerator8x8[1939] = 8'h30;
assign _c_characterGenerator8x8[1940] = 8'h60;
assign _c_characterGenerator8x8[1941] = 8'h00;
assign _c_characterGenerator8x8[1942] = 8'hfc;
assign _c_characterGenerator8x8[1943] = 8'h00;
assign _c_characterGenerator8x8[1944] = 8'h18;
assign _c_characterGenerator8x8[1945] = 8'h30;
assign _c_characterGenerator8x8[1946] = 8'h60;
assign _c_characterGenerator8x8[1947] = 8'h30;
assign _c_characterGenerator8x8[1948] = 8'h18;
assign _c_characterGenerator8x8[1949] = 8'h00;
assign _c_characterGenerator8x8[1950] = 8'hfc;
assign _c_characterGenerator8x8[1951] = 8'h00;
assign _c_characterGenerator8x8[1952] = 8'h0e;
assign _c_characterGenerator8x8[1953] = 8'h1b;
assign _c_characterGenerator8x8[1954] = 8'h1b;
assign _c_characterGenerator8x8[1955] = 8'h18;
assign _c_characterGenerator8x8[1956] = 8'h18;
assign _c_characterGenerator8x8[1957] = 8'h18;
assign _c_characterGenerator8x8[1958] = 8'h18;
assign _c_characterGenerator8x8[1959] = 8'h18;
assign _c_characterGenerator8x8[1960] = 8'h18;
assign _c_characterGenerator8x8[1961] = 8'h18;
assign _c_characterGenerator8x8[1962] = 8'h18;
assign _c_characterGenerator8x8[1963] = 8'h18;
assign _c_characterGenerator8x8[1964] = 8'h18;
assign _c_characterGenerator8x8[1965] = 8'hd8;
assign _c_characterGenerator8x8[1966] = 8'hd8;
assign _c_characterGenerator8x8[1967] = 8'h70;
assign _c_characterGenerator8x8[1968] = 8'h30;
assign _c_characterGenerator8x8[1969] = 8'h30;
assign _c_characterGenerator8x8[1970] = 8'h00;
assign _c_characterGenerator8x8[1971] = 8'hfc;
assign _c_characterGenerator8x8[1972] = 8'h00;
assign _c_characterGenerator8x8[1973] = 8'h30;
assign _c_characterGenerator8x8[1974] = 8'h30;
assign _c_characterGenerator8x8[1975] = 8'h00;
assign _c_characterGenerator8x8[1976] = 8'h00;
assign _c_characterGenerator8x8[1977] = 8'h76;
assign _c_characterGenerator8x8[1978] = 8'hdc;
assign _c_characterGenerator8x8[1979] = 8'h00;
assign _c_characterGenerator8x8[1980] = 8'h76;
assign _c_characterGenerator8x8[1981] = 8'hdc;
assign _c_characterGenerator8x8[1982] = 8'h00;
assign _c_characterGenerator8x8[1983] = 8'h00;
assign _c_characterGenerator8x8[1984] = 8'h38;
assign _c_characterGenerator8x8[1985] = 8'h6c;
assign _c_characterGenerator8x8[1986] = 8'h6c;
assign _c_characterGenerator8x8[1987] = 8'h38;
assign _c_characterGenerator8x8[1988] = 8'h00;
assign _c_characterGenerator8x8[1989] = 8'h00;
assign _c_characterGenerator8x8[1990] = 8'h00;
assign _c_characterGenerator8x8[1991] = 8'h00;
assign _c_characterGenerator8x8[1992] = 8'h00;
assign _c_characterGenerator8x8[1993] = 8'h00;
assign _c_characterGenerator8x8[1994] = 8'h00;
assign _c_characterGenerator8x8[1995] = 8'h18;
assign _c_characterGenerator8x8[1996] = 8'h18;
assign _c_characterGenerator8x8[1997] = 8'h00;
assign _c_characterGenerator8x8[1998] = 8'h00;
assign _c_characterGenerator8x8[1999] = 8'h00;
assign _c_characterGenerator8x8[2000] = 8'h00;
assign _c_characterGenerator8x8[2001] = 8'h00;
assign _c_characterGenerator8x8[2002] = 8'h00;
assign _c_characterGenerator8x8[2003] = 8'h00;
assign _c_characterGenerator8x8[2004] = 8'h18;
assign _c_characterGenerator8x8[2005] = 8'h00;
assign _c_characterGenerator8x8[2006] = 8'h00;
assign _c_characterGenerator8x8[2007] = 8'h00;
assign _c_characterGenerator8x8[2008] = 8'h0f;
assign _c_characterGenerator8x8[2009] = 8'h0c;
assign _c_characterGenerator8x8[2010] = 8'h0c;
assign _c_characterGenerator8x8[2011] = 8'h0c;
assign _c_characterGenerator8x8[2012] = 8'hec;
assign _c_characterGenerator8x8[2013] = 8'h6c;
assign _c_characterGenerator8x8[2014] = 8'h3c;
assign _c_characterGenerator8x8[2015] = 8'h1c;
assign _c_characterGenerator8x8[2016] = 8'h78;
assign _c_characterGenerator8x8[2017] = 8'h6c;
assign _c_characterGenerator8x8[2018] = 8'h6c;
assign _c_characterGenerator8x8[2019] = 8'h6c;
assign _c_characterGenerator8x8[2020] = 8'h6c;
assign _c_characterGenerator8x8[2021] = 8'h00;
assign _c_characterGenerator8x8[2022] = 8'h00;
assign _c_characterGenerator8x8[2023] = 8'h00;
assign _c_characterGenerator8x8[2024] = 8'h70;
assign _c_characterGenerator8x8[2025] = 8'h18;
assign _c_characterGenerator8x8[2026] = 8'h30;
assign _c_characterGenerator8x8[2027] = 8'h60;
assign _c_characterGenerator8x8[2028] = 8'h78;
assign _c_characterGenerator8x8[2029] = 8'h00;
assign _c_characterGenerator8x8[2030] = 8'h00;
assign _c_characterGenerator8x8[2031] = 8'h00;
assign _c_characterGenerator8x8[2032] = 8'h00;
assign _c_characterGenerator8x8[2033] = 8'h00;
assign _c_characterGenerator8x8[2034] = 8'h3c;
assign _c_characterGenerator8x8[2035] = 8'h3c;
assign _c_characterGenerator8x8[2036] = 8'h3c;
assign _c_characterGenerator8x8[2037] = 8'h3c;
assign _c_characterGenerator8x8[2038] = 8'h00;
assign _c_characterGenerator8x8[2039] = 8'h00;
assign _c_characterGenerator8x8[2040] = 8'h00;
assign _c_characterGenerator8x8[2041] = 8'h00;
assign _c_characterGenerator8x8[2042] = 8'h00;
assign _c_characterGenerator8x8[2043] = 8'h00;
assign _c_characterGenerator8x8[2044] = 8'h00;
assign _c_characterGenerator8x8[2045] = 8'h00;
assign _c_characterGenerator8x8[2046] = 8'h00;
assign _c_characterGenerator8x8[2047] = 8'h00;
wire  [7:0] _c_character_wdata0;
assign _c_character_wdata0 = 0;
wire  [7:0] _c_foreground_wdata0;
assign _c_foreground_wdata0 = 0;
wire  [7:0] _c_background_wdata0;
assign _c_background_wdata0 = 0;
wire  [7:0] _c_terminal_wdata0;
assign _c_terminal_wdata0 = 0;
wire  [7:0] _c_terminal_y;
assign _c_terminal_y = 3;
wire  [7:0] _c_bitmap_wdata0;
assign _c_bitmap_wdata0 = 0;
wire  [5:0] _c_colourexpand3to6[7:0];
assign _c_colourexpand3to6[0] = 0;
assign _c_colourexpand3to6[1] = 9;
assign _c_colourexpand3to6[2] = 18;
assign _c_colourexpand3to6[3] = 27;
assign _c_colourexpand3to6[4] = 36;
assign _c_colourexpand3to6[5] = 45;
assign _c_colourexpand3to6[6] = 54;
assign _c_colourexpand3to6[7] = 63;
wire  [5:0] _c_colourexpand2to6[3:0];
assign _c_colourexpand2to6[0] = 0;
assign _c_colourexpand2to6[1] = 21;
assign _c_colourexpand2to6[2] = 42;
assign _c_colourexpand2to6[3] = 63;
wire signed [15:0] _c_gpu_temp1;
assign _c_gpu_temp1 = 0;
wire  [7:0] _w_xcharacterpos;
wire  [11:0] _w_ycharacterpos;
wire  [7:0] _w_xincharacter;
wire  [7:0] _w_yincharacter;
wire  [0:0] _w_characterpixel;
wire  [7:0] _w_xterminalpos;
wire  [11:0] _w_yterminalpos;
wire  [0:0] _w_is_cursor;
wire  [7:0] _w_xinterminal;
wire  [7:0] _w_yinterminal;
wire  [0:0] _w_terminalpixel;

reg  [0:0] _d_character_wenable0;
reg  [0:0] _q_character_wenable0;
reg  [11:0] _d_character_addr0;
reg  [11:0] _q_character_addr0;
reg  [0:0] _d_character_wenable1;
reg  [0:0] _q_character_wenable1;
reg  [7:0] _d_character_wdata1;
reg  [7:0] _q_character_wdata1;
reg  [11:0] _d_character_addr1;
reg  [11:0] _q_character_addr1;
reg  [0:0] _d_foreground_wenable0;
reg  [0:0] _q_foreground_wenable0;
reg  [11:0] _d_foreground_addr0;
reg  [11:0] _q_foreground_addr0;
reg  [0:0] _d_foreground_wenable1;
reg  [0:0] _q_foreground_wenable1;
reg  [7:0] _d_foreground_wdata1;
reg  [7:0] _q_foreground_wdata1;
reg  [11:0] _d_foreground_addr1;
reg  [11:0] _q_foreground_addr1;
reg  [0:0] _d_background_wenable0;
reg  [0:0] _q_background_wenable0;
reg  [11:0] _d_background_addr0;
reg  [11:0] _q_background_addr0;
reg  [0:0] _d_background_wenable1;
reg  [0:0] _q_background_wenable1;
reg  [7:0] _d_background_wdata1;
reg  [7:0] _q_background_wdata1;
reg  [11:0] _d_background_addr1;
reg  [11:0] _q_background_addr1;
reg  [0:0] _d_terminal_wenable0;
reg  [0:0] _q_terminal_wenable0;
reg  [8:0] _d_terminal_addr0;
reg  [8:0] _q_terminal_addr0;
reg  [0:0] _d_terminal_wenable1;
reg  [0:0] _q_terminal_wenable1;
reg  [7:0] _d_terminal_wdata1;
reg  [7:0] _q_terminal_wdata1;
reg  [8:0] _d_terminal_addr1;
reg  [8:0] _q_terminal_addr1;
reg  [7:0] _d_terminal_x;
reg  [7:0] _q_terminal_x;
reg  [1:0] _d_terminal_active;
reg  [1:0] _q_terminal_active;
reg  [8:0] _d_terminal_scroll;
reg  [8:0] _q_terminal_scroll;
reg  [7:0] _d_terminal_scroll_next;
reg  [7:0] _q_terminal_scroll_next;
reg  [0:0] _d_bitmap_wenable0;
reg  [0:0] _q_bitmap_wenable0;
reg  [18:0] _d_bitmap_addr0;
reg  [18:0] _q_bitmap_addr0;
reg  [0:0] _d_bitmap_wenable1;
reg  [0:0] _q_bitmap_wenable1;
reg  [7:0] _d_bitmap_wdata1;
reg  [7:0] _q_bitmap_wdata1;
reg  [18:0] _d_bitmap_addr1;
reg  [18:0] _q_bitmap_addr1;
reg  [15:0] _d_gpu_active_x;
reg  [15:0] _q_gpu_active_x;
reg  [15:0] _d_gpu_active_y;
reg  [15:0] _q_gpu_active_y;
reg  [7:0] _d_gpu_active_colour;
reg  [7:0] _q_gpu_active_colour;
reg signed [15:0] _d_gpu_temp0;
reg signed [15:0] _q_gpu_temp0;
reg signed [15:0] _d_gpu_temp2;
reg signed [15:0] _q_gpu_temp2;
reg signed [15:0] _d_gpu_temp3;
reg signed [15:0] _q_gpu_temp3;
reg signed [15:0] _d_gpu_temp4;
reg signed [15:0] _q_gpu_temp4;
reg  [5:0] _d_pix_red,_q_pix_red;
reg  [5:0] _d_pix_green,_q_pix_green;
reg  [5:0] _d_pix_blue,_q_pix_blue;
reg  [7:0] _d_gpu_active,_q_gpu_active;
reg  [1:0] _d_index,_q_index;
assign out_pix_red = _d_pix_red;
assign out_pix_green = _d_pix_green;
assign out_pix_blue = _d_pix_blue;
assign out_gpu_active = _q_gpu_active;
assign out_done = (_q_index == 3);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_character_wenable0 <= 0;
_q_character_addr0 <= 0;
_q_character_wenable1 <= 0;
_q_character_wdata1 <= 0;
_q_character_addr1 <= 0;
_q_foreground_wenable0 <= 0;
_q_foreground_addr0 <= 0;
_q_foreground_wenable1 <= 0;
_q_foreground_wdata1 <= 0;
_q_foreground_addr1 <= 0;
_q_background_wenable0 <= 0;
_q_background_addr0 <= 0;
_q_background_wenable1 <= 0;
_q_background_wdata1 <= 0;
_q_background_addr1 <= 0;
_q_terminal_wenable0 <= 0;
_q_terminal_addr0 <= 0;
_q_terminal_wenable1 <= 0;
_q_terminal_wdata1 <= 0;
_q_terminal_addr1 <= 0;
_q_terminal_x <= 0;
_q_terminal_active <= 0;
_q_terminal_scroll <= 0;
_q_terminal_scroll_next <= 0;
_q_bitmap_wenable0 <= 0;
_q_bitmap_addr0 <= 0;
_q_bitmap_wenable1 <= 0;
_q_bitmap_wdata1 <= 0;
_q_bitmap_addr1 <= 0;
_q_gpu_active_x <= 0;
_q_gpu_active_y <= 0;
_q_gpu_active_colour <= 0;
_q_gpu_temp0 <= 0;
_q_gpu_temp2 <= 0;
_q_gpu_temp3 <= 0;
_q_gpu_temp4 <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_character_wenable0 <= _d_character_wenable0;
_q_character_addr0 <= _d_character_addr0;
_q_character_wenable1 <= _d_character_wenable1;
_q_character_wdata1 <= _d_character_wdata1;
_q_character_addr1 <= _d_character_addr1;
_q_foreground_wenable0 <= _d_foreground_wenable0;
_q_foreground_addr0 <= _d_foreground_addr0;
_q_foreground_wenable1 <= _d_foreground_wenable1;
_q_foreground_wdata1 <= _d_foreground_wdata1;
_q_foreground_addr1 <= _d_foreground_addr1;
_q_background_wenable0 <= _d_background_wenable0;
_q_background_addr0 <= _d_background_addr0;
_q_background_wenable1 <= _d_background_wenable1;
_q_background_wdata1 <= _d_background_wdata1;
_q_background_addr1 <= _d_background_addr1;
_q_terminal_wenable0 <= _d_terminal_wenable0;
_q_terminal_addr0 <= _d_terminal_addr0;
_q_terminal_wenable1 <= _d_terminal_wenable1;
_q_terminal_wdata1 <= _d_terminal_wdata1;
_q_terminal_addr1 <= _d_terminal_addr1;
_q_terminal_x <= _d_terminal_x;
_q_terminal_active <= _d_terminal_active;
_q_terminal_scroll <= _d_terminal_scroll;
_q_terminal_scroll_next <= _d_terminal_scroll_next;
_q_bitmap_wenable0 <= _d_bitmap_wenable0;
_q_bitmap_addr0 <= _d_bitmap_addr0;
_q_bitmap_wenable1 <= _d_bitmap_wenable1;
_q_bitmap_wdata1 <= _d_bitmap_wdata1;
_q_bitmap_addr1 <= _d_bitmap_addr1;
_q_gpu_active_x <= _d_gpu_active_x;
_q_gpu_active_y <= _d_gpu_active_y;
_q_gpu_active_colour <= _d_gpu_active_colour;
_q_gpu_temp0 <= _d_gpu_temp0;
_q_gpu_temp2 <= _d_gpu_temp2;
_q_gpu_temp3 <= _d_gpu_temp3;
_q_gpu_temp4 <= _d_gpu_temp4;
_q_index <= _d_index;
  end
_q_pix_red <= _d_pix_red;
_q_pix_green <= _d_pix_green;
_q_pix_blue <= _d_pix_blue;
_q_gpu_active <= _d_gpu_active;
end


M_multiplex_display_mem_character __mem__character(
.clock0(clock),
.clock1(clock),
.in_character_wenable0(_d_character_wenable0),
.in_character_wdata0(_c_character_wdata0),
.in_character_addr0(_d_character_addr0),
.in_character_wenable1(_d_character_wenable1),
.in_character_wdata1(_d_character_wdata1),
.in_character_addr1(_d_character_addr1),
.out_character_rdata0(_w_mem_character_rdata0),
.out_character_rdata1(_w_mem_character_rdata1)
);
M_multiplex_display_mem_foreground __mem__foreground(
.clock0(clock),
.clock1(clock),
.in_foreground_wenable0(_d_foreground_wenable0),
.in_foreground_wdata0(_c_foreground_wdata0),
.in_foreground_addr0(_d_foreground_addr0),
.in_foreground_wenable1(_d_foreground_wenable1),
.in_foreground_wdata1(_d_foreground_wdata1),
.in_foreground_addr1(_d_foreground_addr1),
.out_foreground_rdata0(_w_mem_foreground_rdata0),
.out_foreground_rdata1(_w_mem_foreground_rdata1)
);
M_multiplex_display_mem_background __mem__background(
.clock0(clock),
.clock1(clock),
.in_background_wenable0(_d_background_wenable0),
.in_background_wdata0(_c_background_wdata0),
.in_background_addr0(_d_background_addr0),
.in_background_wenable1(_d_background_wenable1),
.in_background_wdata1(_d_background_wdata1),
.in_background_addr1(_d_background_addr1),
.out_background_rdata0(_w_mem_background_rdata0),
.out_background_rdata1(_w_mem_background_rdata1)
);
M_multiplex_display_mem_terminal __mem__terminal(
.clock0(clock),
.clock1(clock),
.in_terminal_wenable0(_d_terminal_wenable0),
.in_terminal_wdata0(_c_terminal_wdata0),
.in_terminal_addr0(_d_terminal_addr0),
.in_terminal_wenable1(_d_terminal_wenable1),
.in_terminal_wdata1(_d_terminal_wdata1),
.in_terminal_addr1(_d_terminal_addr1),
.out_terminal_rdata0(_w_mem_terminal_rdata0),
.out_terminal_rdata1(_w_mem_terminal_rdata1)
);
M_multiplex_display_mem_bitmap __mem__bitmap(
.clock0(clock),
.clock1(clock),
.in_bitmap_wenable0(_d_bitmap_wenable0),
.in_bitmap_wdata0(_c_bitmap_wdata0),
.in_bitmap_addr0(_d_bitmap_addr0),
.in_bitmap_wenable1(_d_bitmap_wenable1),
.in_bitmap_wdata1(_d_bitmap_wdata1),
.in_bitmap_addr1(_d_bitmap_addr1),
.out_bitmap_rdata0(_w_mem_bitmap_rdata0),
.out_bitmap_rdata1(_w_mem_bitmap_rdata1)
);

assign _w_terminalpixel = ((_c_characterGenerator8x8[_w_mem_terminal_rdata0*8+_w_yinterminal]<<_w_xinterminal)>>7)&1;
assign _w_yinterminal = in_pix_y&7;
assign _w_xinterminal = in_pix_x&7;
assign _w_is_cursor = (_w_xterminalpos==_d_terminal_x)&(((in_pix_y-448)>>3)==_c_terminal_y);
assign _w_yterminalpos = ((in_pix_y-448)>>3)*80;
assign _w_characterpixel = ((_c_characterGenerator8x16[_w_mem_character_rdata0*16+_w_yincharacter]<<_w_xincharacter)>>7)&1;
assign _w_yincharacter = in_pix_y&15;
assign _w_ycharacterpos = ((in_pix_y)>>4)*80;
assign _w_xterminalpos = (in_pix_x+1)>>3;
assign _w_xincharacter = in_pix_x&7;
assign _w_xcharacterpos = (in_pix_x+1)>>3;

always @* begin
_d_character_wenable0 = _q_character_wenable0;
_d_character_addr0 = _q_character_addr0;
_d_character_wenable1 = _q_character_wenable1;
_d_character_wdata1 = _q_character_wdata1;
_d_character_addr1 = _q_character_addr1;
_d_foreground_wenable0 = _q_foreground_wenable0;
_d_foreground_addr0 = _q_foreground_addr0;
_d_foreground_wenable1 = _q_foreground_wenable1;
_d_foreground_wdata1 = _q_foreground_wdata1;
_d_foreground_addr1 = _q_foreground_addr1;
_d_background_wenable0 = _q_background_wenable0;
_d_background_addr0 = _q_background_addr0;
_d_background_wenable1 = _q_background_wenable1;
_d_background_wdata1 = _q_background_wdata1;
_d_background_addr1 = _q_background_addr1;
_d_terminal_wenable0 = _q_terminal_wenable0;
_d_terminal_addr0 = _q_terminal_addr0;
_d_terminal_wenable1 = _q_terminal_wenable1;
_d_terminal_wdata1 = _q_terminal_wdata1;
_d_terminal_addr1 = _q_terminal_addr1;
_d_terminal_x = _q_terminal_x;
_d_terminal_active = _q_terminal_active;
_d_terminal_scroll = _q_terminal_scroll;
_d_terminal_scroll_next = _q_terminal_scroll_next;
_d_bitmap_wenable0 = _q_bitmap_wenable0;
_d_bitmap_addr0 = _q_bitmap_addr0;
_d_bitmap_wenable1 = _q_bitmap_wenable1;
_d_bitmap_wdata1 = _q_bitmap_wdata1;
_d_bitmap_addr1 = _q_bitmap_addr1;
_d_gpu_active_x = _q_gpu_active_x;
_d_gpu_active_y = _q_gpu_active_y;
_d_gpu_active_colour = _q_gpu_active_colour;
_d_gpu_temp0 = _q_gpu_temp0;
_d_gpu_temp2 = _q_gpu_temp2;
_d_gpu_temp3 = _q_gpu_temp3;
_d_gpu_temp4 = _q_gpu_temp4;
_d_pix_red = _q_pix_red;
_d_pix_green = _q_pix_green;
_d_pix_blue = _q_pix_blue;
_d_gpu_active = _q_gpu_active;
_d_index = _q_index;
// _always_pre
_d_pix_red = 0;
_d_pix_green = 0;
_d_pix_blue = 0;
_d_terminal_addr0 = _w_xterminalpos+_w_yterminalpos;
_d_terminal_wenable0 = 0;
_d_character_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_character_wenable0 = 0;
_d_foreground_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_foreground_wenable0 = 0;
_d_background_addr0 = _w_xcharacterpos+_w_ycharacterpos;
_d_background_wenable0 = 0;
_d_bitmap_addr0 = in_pix_x+in_pix_y*640;
_d_bitmap_wenable0 = 0;
_d_bitmap_wenable1 = 0;
_d_character_addr1 = in_tpu_x+in_tpu_y*80;
_d_character_wenable1 = 0;
_d_background_addr1 = in_tpu_x+in_tpu_y*80;
_d_background_wenable1 = 0;
_d_foreground_addr1 = in_tpu_x+in_tpu_y*80;
_d_foreground_wenable1 = 0;
_d_terminal_wenable1 = 0;
_d_index = 3;
case (_q_index)
0: begin
// _top
// var inits
_d_character_wenable0 = 0;
_d_character_addr0 = 0;
_d_character_wenable1 = 0;
_d_character_wdata1 = 0;
_d_character_addr1 = 0;
_d_foreground_wenable0 = 0;
_d_foreground_addr0 = 0;
_d_foreground_wenable1 = 0;
_d_foreground_wdata1 = 0;
_d_foreground_addr1 = 0;
_d_background_wenable0 = 0;
_d_background_addr0 = 0;
_d_background_wenable1 = 0;
_d_background_wdata1 = 0;
_d_background_addr1 = 0;
_d_terminal_wenable0 = 0;
_d_terminal_addr0 = 0;
_d_terminal_wenable1 = 0;
_d_terminal_wdata1 = 0;
_d_terminal_addr1 = 0;
_d_terminal_x = 0;
_d_terminal_active = 0;
_d_terminal_scroll = 0;
_d_terminal_scroll_next = 0;
_d_bitmap_wenable0 = 0;
_d_bitmap_addr0 = 0;
_d_bitmap_wenable1 = 0;
_d_bitmap_wdata1 = 0;
_d_bitmap_addr1 = 0;
_d_gpu_active_x = 0;
_d_gpu_active_y = 0;
_d_gpu_active_colour = 0;
_d_gpu_temp0 = 0;
_d_gpu_temp2 = 0;
_d_gpu_temp3 = 0;
_d_gpu_temp4 = 0;
// --
_d_gpu_active = 0;
_d_index = 1;
end
1: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
  case (in_tpu_write)
  1: begin
// __block_6_case
// __block_7
_d_character_wdata1 = in_tpu_set;
_d_character_wenable1 = 1;
// __block_8
  end
  2: begin
// __block_9_case
// __block_10
_d_background_wdata1 = in_tpu_set;
_d_background_wenable1 = 1;
// __block_11
  end
  3: begin
// __block_12_case
// __block_13
_d_foreground_wdata1 = in_tpu_set;
_d_foreground_wenable1 = 1;
// __block_14
  end
  default: begin
// __block_15_case
// __block_16
// __block_17
  end
endcase
// __block_5
if (_q_terminal_active==0) begin
// __block_18
// __block_20
  case (in_terminal_write)
  1: begin
// __block_22_case
// __block_23
  case (in_terminal_character)
  10: begin
// __block_25_case
// __block_26
_d_terminal_scroll = 0;
_d_terminal_active = 1;
// __block_27
  end
  13: begin
// __block_28_case
// __block_29
_d_terminal_x = 0;
_d_terminal_active = 1;
// __block_30
  end
  default: begin
// __block_31_case
// __block_32
_d_terminal_addr1 = _q_terminal_x+_c_terminal_y*80;
_d_terminal_wdata1 = in_terminal_character;
_d_terminal_wenable1 = 1;
if (_q_terminal_x==79) begin
// __block_33
// __block_35
_d_terminal_x = 0;
_d_terminal_scroll = 0;
_d_terminal_active = 1;
// __block_36
end else begin
// __block_34
// __block_37
_d_terminal_x = _q_terminal_x+1;
// __block_38
end
// __block_39
// __block_40
  end
endcase
// __block_24
// __block_41
  end
  default: begin
// __block_42_case
// __block_43
// __block_44
  end
endcase
// __block_21
// __block_45
end else begin
// __block_19
// __block_46
  case (_q_terminal_active)
  1: begin
// __block_48_case
// __block_49
if (_q_terminal_scroll==240) begin
// __block_50
// __block_52
_d_terminal_active = 4;
// __block_53
end else begin
// __block_51
// __block_54
_d_terminal_addr1 = _q_terminal_scroll+80;
_d_terminal_active = 2;
// __block_55
end
// __block_56
// __block_57
  end
  2: begin
// __block_58_case
// __block_59
_d_terminal_scroll_next = _w_mem_terminal_rdata1;
_d_terminal_active = 3;
// __block_60
  end
  3: begin
// __block_61_case
// __block_62
_d_terminal_addr1 = _q_terminal_scroll;
_d_terminal_wdata1 = _q_terminal_scroll_next;
_d_terminal_wenable1 = 1;
_d_terminal_scroll = _q_terminal_scroll+1;
_d_terminal_active = 1;
// __block_63
  end
  4: begin
// __block_64_case
// __block_65
_d_terminal_addr1 = _q_terminal_scroll;
_d_terminal_wdata1 = 0;
_d_terminal_wenable1 = 1;
if (_q_terminal_scroll==320) begin
// __block_66
// __block_68
_d_terminal_active = 0;
// __block_69
end else begin
// __block_67
// __block_70
_d_terminal_scroll = _q_terminal_scroll+1;
// __block_71
end
// __block_72
// __block_73
  end
  default: begin
// __block_74_case
// __block_75
// __block_76
  end
endcase
// __block_47
// __block_77
end
// __block_78
  case (_q_gpu_active)
  0: begin
// __block_80_case
// __block_81
  case (in_gpu_write)
  1: begin
// __block_83_case
// __block_84
_d_gpu_active_colour = in_gpu_colour;
_d_gpu_active_x = in_gpu_x;
_d_gpu_active_y = in_gpu_y;
_d_gpu_active = 1;
// __block_85
  end
  2: begin
// __block_86_case
// __block_87
_d_gpu_active_colour = in_gpu_colour;
_d_gpu_active_x = (in_gpu_x<in_gpu_param0)?in_gpu_x:in_gpu_param0;
_d_gpu_active_y = (in_gpu_y<in_gpu_param1)?in_gpu_y:in_gpu_param1;
_d_gpu_temp0 = (in_gpu_x<in_gpu_param0)?in_gpu_x:in_gpu_param0;
_d_gpu_temp2 = (in_gpu_x<in_gpu_param0)?in_gpu_param0:in_gpu_x;
_d_gpu_temp3 = (in_gpu_y<in_gpu_param1)?in_gpu_param1:in_gpu_y;
_d_gpu_active = 2;
// __block_88
  end
  3: begin
// __block_89_case
// __block_90
_d_gpu_active_colour = in_gpu_colour;
_d_gpu_active_x = in_gpu_x;
_d_gpu_active_y = in_gpu_y;
_d_gpu_temp0 = in_gpu_param0;
_d_gpu_temp2 = in_gpu_param0-in_gpu_x;
_d_gpu_temp3 = in_gpu_param1-in_gpu_y;
if ((in_gpu_param0-in_gpu_x)>=(in_gpu_param1-in_gpu_y)) begin
// __block_91
// __block_93
_d_gpu_temp4 = 2*((in_gpu_param1-in_gpu_y)-(in_gpu_param0-in_gpu_x));
_d_gpu_active = 3;
// __block_94
end else begin
// __block_92
// __block_95
_d_gpu_temp4 = 2*((in_gpu_param1-in_gpu_y)-(in_gpu_param0-in_gpu_x));
_d_gpu_active = 4;
// __block_96
end
// __block_97
// __block_98
  end
  default: begin
// __block_99_case
// __block_100
// __block_101
  end
endcase
// __block_82
// __block_102
  end
  1: begin
// __block_103_case
// __block_104
_d_bitmap_addr1 = _q_gpu_active_x+_q_gpu_active_y*640;
_d_bitmap_wdata1 = _q_gpu_active_colour;
_d_bitmap_wenable1 = 1;
_d_gpu_active = 0;
// __block_105
  end
  2: begin
// __block_106_case
// __block_107
_d_bitmap_addr1 = _q_gpu_active_x+_q_gpu_active_y*640;
_d_bitmap_wdata1 = _q_gpu_active_colour;
_d_bitmap_wenable1 = 1;
if (_q_gpu_active_x==_q_gpu_temp2) begin
// __block_108
// __block_110
if (_q_gpu_active_y==_q_gpu_temp3) begin
// __block_111
// __block_113
_d_gpu_active = 0;
// __block_114
end else begin
// __block_112
// __block_115
_d_gpu_active_x = _q_gpu_temp0;
_d_gpu_active_y = _q_gpu_active_y+1;
// __block_116
end
// __block_117
// __block_118
end else begin
// __block_109
// __block_119
_d_gpu_active_x = _q_gpu_active_x+1;
// __block_120
end
// __block_121
// __block_122
  end
  3: begin
// __block_123_case
// __block_124
if (_q_gpu_active_x<_q_gpu_temp0) begin
// __block_125
// __block_127
_d_bitmap_addr1 = _q_gpu_active_x+_q_gpu_active_y*640;
_d_bitmap_wdata1 = _q_gpu_active_colour;
_d_bitmap_wenable1 = 1;
if (_q_gpu_temp4>=0) begin
// __block_128
// __block_130
_d_gpu_active_y = _q_gpu_active_y+1;
_d_gpu_temp4 = _q_gpu_temp4+2*_q_gpu_temp3-2*_q_gpu_temp2;
// __block_131
end else begin
// __block_129
// __block_132
_d_gpu_temp4 = _q_gpu_temp4+2*_q_gpu_temp3;
// __block_133
end
// __block_134
_d_gpu_active_x = _q_gpu_active_x+1;
// __block_135
end else begin
// __block_126
// __block_136
_d_gpu_active = 0;
// __block_137
end
// __block_138
// __block_139
  end
  4: begin
// __block_140_case
// __block_141
if (_q_gpu_active_y<_c_gpu_temp1) begin
// __block_142
// __block_144
_d_bitmap_addr1 = _q_gpu_active_x+_q_gpu_active_y*640;
_d_bitmap_wdata1 = _q_gpu_active_colour;
_d_bitmap_wenable1 = 1;
if (_q_gpu_temp4>=0) begin
// __block_145
// __block_147
_d_gpu_active_x = _q_gpu_active_x+1;
_d_gpu_temp4 = _q_gpu_temp4+2*_q_gpu_temp3-2*_q_gpu_temp2;
// __block_148
end else begin
// __block_146
// __block_149
_d_gpu_temp4 = _q_gpu_temp4+2*_q_gpu_temp3;
// __block_150
end
// __block_151
_d_gpu_active_y = _q_gpu_active_y+1;
// __block_152
end else begin
// __block_143
// __block_153
_d_gpu_active = 0;
// __block_154
end
// __block_155
// __block_156
  end
  default: begin
// __block_157_case
// __block_158
_d_gpu_active = 0;
// __block_159
  end
endcase
// __block_79
if (in_pix_vblank==0) begin
// __block_160
// __block_162
if (in_pix_active) begin
// __block_163
// __block_165
if (in_pix_y>447&in_showterminal) begin
// __block_166
// __block_168
  case (_w_terminalpixel)
  0: begin
// __block_170_case
// __block_171
if (_w_is_cursor&in_timer1hz) begin
// __block_172
// __block_174
_d_pix_red = 63;
_d_pix_green = 63;
_d_pix_blue = 63;
// __block_175
end else begin
// __block_173
// __block_176
_d_pix_red = 0;
_d_pix_green = 0;
_d_pix_blue = 63;
// __block_177
end
// __block_178
// __block_179
  end
  1: begin
// __block_180_case
// __block_181
if (_w_is_cursor&in_timer1hz) begin
// __block_182
// __block_184
_d_pix_red = 0;
_d_pix_green = 0;
_d_pix_blue = 63;
// __block_185
end else begin
// __block_183
// __block_186
_d_pix_red = 63;
_d_pix_green = 63;
_d_pix_blue = 63;
// __block_187
end
// __block_188
// __block_189
  end
endcase
// __block_169
// __block_190
end else begin
// __block_167
// __block_191
  case (_w_mem_character_rdata0)
  0: begin
// __block_193_case
// __block_194
_d_pix_red = _c_colourexpand3to6[(_w_mem_bitmap_rdata0&8'he0)>>5];
_d_pix_green = _c_colourexpand3to6[(_w_mem_bitmap_rdata0&8'h1c)>>2];
_d_pix_blue = _c_colourexpand2to6[(_w_mem_bitmap_rdata0&8'h3)];
// __block_195
  end
  default: begin
// __block_196_case
// __block_197
  case (_w_characterpixel)
  0: begin
// __block_199_case
// __block_200
_d_pix_red = _c_colourexpand3to6[(_w_mem_background_rdata0&8'he0)>>5];
_d_pix_green = _c_colourexpand3to6[(_w_mem_background_rdata0&8'h1c)>>2];
_d_pix_blue = _c_colourexpand2to6[(_w_mem_background_rdata0&8'h3)];
// __block_201
  end
  1: begin
// __block_202_case
// __block_203
_d_pix_red = _c_colourexpand3to6[(_w_mem_foreground_rdata0&8'he0)>>5];
_d_pix_green = _c_colourexpand3to6[(_w_mem_foreground_rdata0&8'h1c)>>2];
_d_pix_blue = _c_colourexpand2to6[(_w_mem_foreground_rdata0&8'h3)];
// __block_204
  end
endcase
// __block_198
// __block_205
  end
endcase
// __block_192
// __block_206
end
// __block_207
// __block_208
end else begin
// __block_164
end
// __block_209
// __block_210
end else begin
// __block_161
end
// __block_211
// __block_212
_d_index = 1;
end else begin
_d_index = 2;
end
end
2: begin
// __block_3
_d_index = 3;
end
3: begin // end of multiplex_display
end
default: begin 
_d_index = 3;
 end
endcase
end
endmodule


module M_main_mem_dstack(
input                  [0:0] in_dstack_wenable,
input       [15:0]    in_dstack_wdata,
input                  [7:0]    in_dstack_addr,
output reg  [15:0]    out_dstack_rdata,
input                                      clock
);
reg  [15:0] buffer[255:0];
always @(posedge clock) begin
  if (in_dstack_wenable) begin
    buffer[in_dstack_addr] <= in_dstack_wdata;
  end
  out_dstack_rdata <= buffer[in_dstack_addr];
end

endmodule

module M_main_mem_rstack(
input                  [0:0] in_rstack_wenable,
input       [15:0]    in_rstack_wdata,
input                  [7:0]    in_rstack_addr,
output reg  [15:0]    out_rstack_rdata,
input                                      clock
);
reg  [15:0] buffer[255:0];
always @(posedge clock) begin
  if (in_rstack_wenable) begin
    buffer[in_rstack_addr] <= in_rstack_wdata;
  end
  out_rstack_rdata <= buffer[in_rstack_addr];
end

endmodule

module M_main_mem_rom(
input                  [11:0] in_rom_addr,
output reg  [15:0] out_rom_rdata,
input                                   clock
);
reg  [15:0] buffer[3614:0];
always @(posedge clock) begin
   out_rom_rdata <= buffer[in_rom_addr];
end
initial begin
 buffer[0] = 16'h0E07;
 buffer[1] = 16'h0010;
 buffer[2] = 16'h0000;
 buffer[3] = 16'h0000;
 buffer[4] = 16'h0000;
 buffer[5] = 16'h7F00;
 buffer[6] = 16'h1062;
 buffer[7] = 16'h1140;
 buffer[8] = 16'h0000;
 buffer[9] = 16'h0000;
 buffer[10] = 16'h0000;
 buffer[11] = 16'h0000;
 buffer[12] = 16'h0000;
 buffer[13] = 16'h0000;
 buffer[14] = 16'h0000;
 buffer[15] = 16'h0000;
 buffer[16] = 16'h0000;
 buffer[17] = 16'h0000;
 buffer[18] = 16'h0000;
 buffer[19] = 16'h0000;
 buffer[20] = 16'h0000;
 buffer[21] = 16'h0000;
 buffer[22] = 16'h0000;
 buffer[23] = 16'h1C3E;
 buffer[24] = 16'h1C08;
 buffer[25] = 16'h0952;
 buffer[26] = 16'h0964;
 buffer[27] = 16'h1BD4;
 buffer[28] = 16'h0E1E;
 buffer[29] = 16'h0F0A;
 buffer[30] = 16'h1616;
 buffer[31] = 16'h1698;
 buffer[32] = 16'h16C0;
 buffer[33] = 16'h172C;
 buffer[34] = 16'h0000;
 buffer[35] = 16'h0000;
 buffer[36] = 16'h0000;
 buffer[37] = 16'h0000;
 buffer[38] = 16'h0000;
 buffer[39] = 16'h0000;
 buffer[40] = 16'h0000;
 buffer[41] = 16'h0000;
 buffer[42] = 16'h0000;
 buffer[43] = 16'h0000;
 buffer[44] = 16'h0000;
 buffer[45] = 16'h0000;
 buffer[46] = 16'h0000;
 buffer[47] = 16'h0000;
 buffer[48] = 16'h0000;
 buffer[49] = 16'h0000;
 buffer[50] = 16'h0000;
 buffer[51] = 16'h0000;
 buffer[52] = 16'h0000;
 buffer[53] = 16'h0000;
 buffer[54] = 16'h0000;
 buffer[55] = 16'h0000;
 buffer[56] = 16'h0000;
 buffer[57] = 16'h0000;
 buffer[58] = 16'h0000;
 buffer[59] = 16'h0000;
 buffer[60] = 16'h0000;
 buffer[61] = 16'h0000;
 buffer[62] = 16'h0000;
 buffer[63] = 16'h0000;
 buffer[64] = 16'h6003;
 buffer[65] = 16'h6003;
 buffer[66] = 16'h6003;
 buffer[67] = 16'h6003;
 buffer[68] = 16'h6003;
 buffer[69] = 16'h6003;
 buffer[70] = 16'h6003;
 buffer[71] = 16'h6003;
 buffer[72] = 16'h6003;
 buffer[73] = 16'h6003;
 buffer[74] = 16'h6003;
 buffer[75] = 16'h6003;
 buffer[76] = 16'h6003;
 buffer[77] = 16'h6003;
 buffer[78] = 16'h6003;
 buffer[79] = 16'h710C;
 buffer[80] = 16'h6001;
 buffer[81] = 16'h6001;
 buffer[82] = 16'h6001;
 buffer[83] = 16'h6001;
 buffer[84] = 16'h6001;
 buffer[85] = 16'h6001;
 buffer[86] = 16'h6001;
 buffer[87] = 16'h6001;
 buffer[88] = 16'h6001;
 buffer[89] = 16'h6001;
 buffer[90] = 16'h6001;
 buffer[91] = 16'h6001;
 buffer[92] = 16'h6001;
 buffer[93] = 16'h6001;
 buffer[94] = 16'h6001;
 buffer[95] = 16'h700C;
 buffer[96] = 16'h6100;
 buffer[97] = 16'h700C;
 buffer[98] = 16'h404E;
 buffer[99] = 16'h005E;
 buffer[100] = 16'h404D;
 buffer[101] = 16'h005D;
 buffer[102] = 16'h404C;
 buffer[103] = 16'h005C;
 buffer[104] = 16'h404B;
 buffer[105] = 16'h005B;
 buffer[106] = 16'h404A;
 buffer[107] = 16'h005A;
 buffer[108] = 16'h4049;
 buffer[109] = 16'h0059;
 buffer[110] = 16'h4048;
 buffer[111] = 16'h0058;
 buffer[112] = 16'h4047;
 buffer[113] = 16'h0057;
 buffer[114] = 16'h4046;
 buffer[115] = 16'h0056;
 buffer[116] = 16'h4045;
 buffer[117] = 16'h0055;
 buffer[118] = 16'h4044;
 buffer[119] = 16'h0054;
 buffer[120] = 16'h4043;
 buffer[121] = 16'h0053;
 buffer[122] = 16'h4042;
 buffer[123] = 16'h0052;
 buffer[124] = 16'h4041;
 buffer[125] = 16'h0051;
 buffer[126] = 16'h4040;
 buffer[127] = 16'h0050;
 buffer[128] = 16'h700C;
 buffer[129] = 16'h0000;
 buffer[130] = 16'h0000;
 buffer[131] = 16'h0000;
 buffer[132] = 16'h0000;
 buffer[133] = 16'h0000;
 buffer[134] = 16'h0000;
 buffer[135] = 16'h0000;
 buffer[136] = 16'h0000;
 buffer[137] = 16'h0000;
 buffer[138] = 16'h0000;
 buffer[139] = 16'h0000;
 buffer[140] = 16'h0000;
 buffer[141] = 16'h0000;
 buffer[142] = 16'h0000;
 buffer[143] = 16'h0000;
 buffer[144] = 16'h0000;
 buffer[145] = 16'h0000;
 buffer[146] = 16'h0000;
 buffer[147] = 16'h0000;
 buffer[148] = 16'h0000;
 buffer[149] = 16'h0000;
 buffer[150] = 16'h0000;
 buffer[151] = 16'h0000;
 buffer[152] = 16'h0000;
 buffer[153] = 16'h0000;
 buffer[154] = 16'h0000;
 buffer[155] = 16'h0000;
 buffer[156] = 16'h0000;
 buffer[157] = 16'h0000;
 buffer[158] = 16'h0000;
 buffer[159] = 16'h0000;
 buffer[160] = 16'h0000;
 buffer[161] = 16'h0000;
 buffer[162] = 16'h0000;
 buffer[163] = 16'h0000;
 buffer[164] = 16'h0000;
 buffer[165] = 16'h0000;
 buffer[166] = 16'h0000;
 buffer[167] = 16'h0000;
 buffer[168] = 16'h0000;
 buffer[169] = 16'h0000;
 buffer[170] = 16'h0000;
 buffer[171] = 16'h0000;
 buffer[172] = 16'h0000;
 buffer[173] = 16'h0000;
 buffer[174] = 16'h0000;
 buffer[175] = 16'h0000;
 buffer[176] = 16'h0000;
 buffer[177] = 16'h0000;
 buffer[178] = 16'h0000;
 buffer[179] = 16'h0000;
 buffer[180] = 16'h0000;
 buffer[181] = 16'h0000;
 buffer[182] = 16'h0000;
 buffer[183] = 16'h0000;
 buffer[184] = 16'h0000;
 buffer[185] = 16'h0000;
 buffer[186] = 16'h0000;
 buffer[187] = 16'h0000;
 buffer[188] = 16'h0000;
 buffer[189] = 16'h0000;
 buffer[190] = 16'h0000;
 buffer[191] = 16'h0000;
 buffer[192] = 16'h0000;
 buffer[193] = 16'h6E04;
 buffer[194] = 16'h6F6F;
 buffer[195] = 16'h0070;
 buffer[196] = 16'h700C;
 buffer[197] = 16'h0182;
 buffer[198] = 16'h2B01;
 buffer[199] = 16'h720F;
 buffer[200] = 16'h018C;
 buffer[201] = 16'h7803;
 buffer[202] = 16'h726F;
 buffer[203] = 16'h750F;
 buffer[204] = 16'h0192;
 buffer[205] = 16'h6103;
 buffer[206] = 16'h646E;
 buffer[207] = 16'h730F;
 buffer[208] = 16'h019A;
 buffer[209] = 16'h6F02;
 buffer[210] = 16'h0072;
 buffer[211] = 16'h740F;
 buffer[212] = 16'h01A2;
 buffer[213] = 16'h6906;
 buffer[214] = 16'h766E;
 buffer[215] = 16'h7265;
 buffer[216] = 16'h0074;
 buffer[217] = 16'h760C;
 buffer[218] = 16'h01AA;
 buffer[219] = 16'h3D01;
 buffer[220] = 16'h770F;
 buffer[221] = 16'h01B6;
 buffer[222] = 16'h3C01;
 buffer[223] = 16'h780F;
 buffer[224] = 16'h01BC;
 buffer[225] = 16'h7502;
 buffer[226] = 16'h003C;
 buffer[227] = 16'h7F0F;
 buffer[228] = 16'h01C2;
 buffer[229] = 16'h7304;
 buffer[230] = 16'h6177;
 buffer[231] = 16'h0070;
 buffer[232] = 16'h718C;
 buffer[233] = 16'h01CA;
 buffer[234] = 16'h7502;
 buffer[235] = 16'h003E;
 buffer[236] = 16'h771F;
 buffer[237] = 16'h01D4;
 buffer[238] = 16'h6403;
 buffer[239] = 16'h7075;
 buffer[240] = 16'h708D;
 buffer[241] = 16'h01DC;
 buffer[242] = 16'h6404;
 buffer[243] = 16'h6F72;
 buffer[244] = 16'h0070;
 buffer[245] = 16'h710F;
 buffer[246] = 16'h01E4;
 buffer[247] = 16'h6F04;
 buffer[248] = 16'h6576;
 buffer[249] = 16'h0072;
 buffer[250] = 16'h718D;
 buffer[251] = 16'h01EE;
 buffer[252] = 16'h6E03;
 buffer[253] = 16'h7069;
 buffer[254] = 16'h700F;
 buffer[255] = 16'h01F8;
 buffer[256] = 16'h6C06;
 buffer[257] = 16'h6873;
 buffer[258] = 16'h6669;
 buffer[259] = 16'h0074;
 buffer[260] = 16'h7D0F;
 buffer[261] = 16'h0200;
 buffer[262] = 16'h7206;
 buffer[263] = 16'h6873;
 buffer[264] = 16'h6669;
 buffer[265] = 16'h0074;
 buffer[266] = 16'h790F;
 buffer[267] = 16'h020C;
 buffer[268] = 16'h3102;
 buffer[269] = 16'h002D;
 buffer[270] = 16'h7A0C;
 buffer[271] = 16'h0218;
 buffer[272] = 16'h3E42;
 buffer[273] = 16'h0072;
 buffer[274] = 16'h6B8D;
 buffer[275] = 16'h6180;
 buffer[276] = 16'h6147;
 buffer[277] = 16'h6147;
 buffer[278] = 16'h700C;
 buffer[279] = 16'h0220;
 buffer[280] = 16'h7242;
 buffer[281] = 16'h003E;
 buffer[282] = 16'h6B8D;
 buffer[283] = 16'h6B8D;
 buffer[284] = 16'h6180;
 buffer[285] = 16'h6147;
 buffer[286] = 16'h700C;
 buffer[287] = 16'h0230;
 buffer[288] = 16'h7242;
 buffer[289] = 16'h0040;
 buffer[290] = 16'h6B8D;
 buffer[291] = 16'h6B8D;
 buffer[292] = 16'h6081;
 buffer[293] = 16'h6147;
 buffer[294] = 16'h6180;
 buffer[295] = 16'h6147;
 buffer[296] = 16'h700C;
 buffer[297] = 16'h0240;
 buffer[298] = 16'h4001;
 buffer[299] = 16'h7C0C;
 buffer[300] = 16'h0254;
 buffer[301] = 16'h2101;
 buffer[302] = 16'h6023;
 buffer[303] = 16'h710F;
 buffer[304] = 16'h025A;
 buffer[305] = 16'h3C02;
 buffer[306] = 16'h003E;
 buffer[307] = 16'h721F;
 buffer[308] = 16'h0262;
 buffer[309] = 16'h3002;
 buffer[310] = 16'h003C;
 buffer[311] = 16'h781C;
 buffer[312] = 16'h026A;
 buffer[313] = 16'h3002;
 buffer[314] = 16'h003D;
 buffer[315] = 16'h701C;
 buffer[316] = 16'h0272;
 buffer[317] = 16'h3003;
 buffer[318] = 16'h3E3C;
 buffer[319] = 16'h711C;
 buffer[320] = 16'h027A;
 buffer[321] = 16'h3E01;
 buffer[322] = 16'h761F;
 buffer[323] = 16'h0282;
 buffer[324] = 16'h3002;
 buffer[325] = 16'h003E;
 buffer[326] = 16'h791C;
 buffer[327] = 16'h0288;
 buffer[328] = 16'h3E02;
 buffer[329] = 16'h003D;
 buffer[330] = 16'h7F1F;
 buffer[331] = 16'h0290;
 buffer[332] = 16'h7404;
 buffer[333] = 16'h6375;
 buffer[334] = 16'h006B;
 buffer[335] = 16'h6180;
 buffer[336] = 16'h718D;
 buffer[337] = 16'h0298;
 buffer[338] = 16'h2D04;
 buffer[339] = 16'h6F72;
 buffer[340] = 16'h0074;
 buffer[341] = 16'h6180;
 buffer[342] = 16'h6147;
 buffer[343] = 16'h6180;
 buffer[344] = 16'h6B8D;
 buffer[345] = 16'h700C;
 buffer[346] = 16'h02A4;
 buffer[347] = 16'h3202;
 buffer[348] = 16'h002F;
 buffer[349] = 16'h8001;
 buffer[350] = 16'h790F;
 buffer[351] = 16'h02B6;
 buffer[352] = 16'h3202;
 buffer[353] = 16'h002A;
 buffer[354] = 16'h741C;
 buffer[355] = 16'h02C0;
 buffer[356] = 16'h3102;
 buffer[357] = 16'h002B;
 buffer[358] = 16'h731C;
 buffer[359] = 16'h02C8;
 buffer[360] = 16'h7303;
 buffer[361] = 16'h4070;
 buffer[362] = 16'h6E81;
 buffer[363] = 16'h80FF;
 buffer[364] = 16'h730F;
 buffer[365] = 16'h02D0;
 buffer[366] = 16'h6507;
 buffer[367] = 16'h6578;
 buffer[368] = 16'h7563;
 buffer[369] = 16'h6574;
 buffer[370] = 16'h6147;
 buffer[371] = 16'h700C;
 buffer[372] = 16'h02DC;
 buffer[373] = 16'h6203;
 buffer[374] = 16'h6579;
 buffer[375] = 16'h8FFD;
 buffer[376] = 16'h6600;
 buffer[377] = 16'h6023;
 buffer[378] = 16'h710F;
 buffer[379] = 16'h02EA;
 buffer[380] = 16'h6302;
 buffer[381] = 16'h0040;
 buffer[382] = 16'h6081;
 buffer[383] = 16'h6C00;
 buffer[384] = 16'h6180;
 buffer[385] = 16'h8001;
 buffer[386] = 16'h6303;
 buffer[387] = 16'h2187;
 buffer[388] = 16'h8008;
 buffer[389] = 16'h6903;
 buffer[390] = 16'h0189;
 buffer[391] = 16'h80FF;
 buffer[392] = 16'h730F;
 buffer[393] = 16'h700C;
 buffer[394] = 16'h02F8;
 buffer[395] = 16'h6302;
 buffer[396] = 16'h0021;
 buffer[397] = 16'h6180;
 buffer[398] = 16'h80FF;
 buffer[399] = 16'h6303;
 buffer[400] = 16'h6081;
 buffer[401] = 16'h8008;
 buffer[402] = 16'h6D03;
 buffer[403] = 16'h6403;
 buffer[404] = 16'h6180;
 buffer[405] = 16'h414F;
 buffer[406] = 16'h6081;
 buffer[407] = 16'h6C00;
 buffer[408] = 16'h6180;
 buffer[409] = 16'h8001;
 buffer[410] = 16'h6303;
 buffer[411] = 16'h8000;
 buffer[412] = 16'h6703;
 buffer[413] = 16'h80FF;
 buffer[414] = 16'h6503;
 buffer[415] = 16'h6147;
 buffer[416] = 16'h6181;
 buffer[417] = 16'h6503;
 buffer[418] = 16'h6B8D;
 buffer[419] = 16'h6303;
 buffer[420] = 16'h6503;
 buffer[421] = 16'h6180;
 buffer[422] = 16'h6023;
 buffer[423] = 16'h710F;
 buffer[424] = 16'h0316;
 buffer[425] = 16'h7503;
 buffer[426] = 16'h2B6D;
 buffer[427] = 16'h6181;
 buffer[428] = 16'h6181;
 buffer[429] = 16'h6203;
 buffer[430] = 16'h6147;
 buffer[431] = 16'h6B81;
 buffer[432] = 16'h8000;
 buffer[433] = 16'h6F13;
 buffer[434] = 16'h6147;
 buffer[435] = 16'h6181;
 buffer[436] = 16'h6181;
 buffer[437] = 16'h6303;
 buffer[438] = 16'h6810;
 buffer[439] = 16'h6B8D;
 buffer[440] = 16'h6403;
 buffer[441] = 16'h6147;
 buffer[442] = 16'h6403;
 buffer[443] = 16'h6810;
 buffer[444] = 16'h6B8D;
 buffer[445] = 16'h6303;
 buffer[446] = 16'h6600;
 buffer[447] = 16'h6310;
 buffer[448] = 16'h6B8D;
 buffer[449] = 16'h718C;
 buffer[450] = 16'h0352;
 buffer[451] = 16'h6445;
 buffer[452] = 16'h766F;
 buffer[453] = 16'h7261;
 buffer[454] = 16'h6B8D;
 buffer[455] = 16'h700C;
 buffer[456] = 16'h0386;
 buffer[457] = 16'h7502;
 buffer[458] = 16'h0070;
 buffer[459] = 16'h41C6;
 buffer[460] = 16'h7E8C;
 buffer[461] = 16'h0392;
 buffer[462] = 16'h6446;
 buffer[463] = 16'h756F;
 buffer[464] = 16'h6573;
 buffer[465] = 16'h0072;
 buffer[466] = 16'h41CB;
 buffer[467] = 16'h6C00;
 buffer[468] = 16'h6B8D;
 buffer[469] = 16'h6C00;
 buffer[470] = 16'h720F;
 buffer[471] = 16'h039C;
 buffer[472] = 16'h6204;
 buffer[473] = 16'h7361;
 buffer[474] = 16'h0065;
 buffer[475] = 16'hFE80;
 buffer[476] = 16'h700C;
 buffer[477] = 16'h03B0;
 buffer[478] = 16'h7404;
 buffer[479] = 16'h6D65;
 buffer[480] = 16'h0070;
 buffer[481] = 16'hFE82;
 buffer[482] = 16'h700C;
 buffer[483] = 16'h03BC;
 buffer[484] = 16'h3E03;
 buffer[485] = 16'h6E69;
 buffer[486] = 16'hFE84;
 buffer[487] = 16'h700C;
 buffer[488] = 16'h03C8;
 buffer[489] = 16'h2304;
 buffer[490] = 16'h6974;
 buffer[491] = 16'h0062;
 buffer[492] = 16'hFE86;
 buffer[493] = 16'h700C;
 buffer[494] = 16'h03D2;
 buffer[495] = 16'h7403;
 buffer[496] = 16'h6269;
 buffer[497] = 16'hFE88;
 buffer[498] = 16'h700C;
 buffer[499] = 16'h03DE;
 buffer[500] = 16'h2705;
 buffer[501] = 16'h7665;
 buffer[502] = 16'h6C61;
 buffer[503] = 16'hFE8A;
 buffer[504] = 16'h700C;
 buffer[505] = 16'h03E8;
 buffer[506] = 16'h2706;
 buffer[507] = 16'h6261;
 buffer[508] = 16'h726F;
 buffer[509] = 16'h0074;
 buffer[510] = 16'hFE8C;
 buffer[511] = 16'h700C;
 buffer[512] = 16'h03F4;
 buffer[513] = 16'h6803;
 buffer[514] = 16'h646C;
 buffer[515] = 16'hFE8E;
 buffer[516] = 16'h700C;
 buffer[517] = 16'h0402;
 buffer[518] = 16'h6307;
 buffer[519] = 16'h6E6F;
 buffer[520] = 16'h6574;
 buffer[521] = 16'h7478;
 buffer[522] = 16'hFE90;
 buffer[523] = 16'h700C;
 buffer[524] = 16'h040C;
 buffer[525] = 16'h660E;
 buffer[526] = 16'h726F;
 buffer[527] = 16'h6874;
 buffer[528] = 16'h772D;
 buffer[529] = 16'h726F;
 buffer[530] = 16'h6C64;
 buffer[531] = 16'h7369;
 buffer[532] = 16'h0074;
 buffer[533] = 16'hFEA2;
 buffer[534] = 16'h700C;
 buffer[535] = 16'h041A;
 buffer[536] = 16'h6307;
 buffer[537] = 16'h7275;
 buffer[538] = 16'h6572;
 buffer[539] = 16'h746E;
 buffer[540] = 16'hFEA8;
 buffer[541] = 16'h700C;
 buffer[542] = 16'h0430;
 buffer[543] = 16'h6402;
 buffer[544] = 16'h0070;
 buffer[545] = 16'hFEAC;
 buffer[546] = 16'h700C;
 buffer[547] = 16'h043E;
 buffer[548] = 16'h6C04;
 buffer[549] = 16'h7361;
 buffer[550] = 16'h0074;
 buffer[551] = 16'hFEAE;
 buffer[552] = 16'h700C;
 buffer[553] = 16'h0448;
 buffer[554] = 16'h2705;
 buffer[555] = 16'h6B3F;
 buffer[556] = 16'h7965;
 buffer[557] = 16'hFEB0;
 buffer[558] = 16'h700C;
 buffer[559] = 16'h0454;
 buffer[560] = 16'h2705;
 buffer[561] = 16'h6D65;
 buffer[562] = 16'h7469;
 buffer[563] = 16'hFEB2;
 buffer[564] = 16'h700C;
 buffer[565] = 16'h0460;
 buffer[566] = 16'h2705;
 buffer[567] = 16'h6F62;
 buffer[568] = 16'h746F;
 buffer[569] = 16'hFEB4;
 buffer[570] = 16'h700C;
 buffer[571] = 16'h046C;
 buffer[572] = 16'h2702;
 buffer[573] = 16'h005C;
 buffer[574] = 16'hFEB6;
 buffer[575] = 16'h700C;
 buffer[576] = 16'h0478;
 buffer[577] = 16'h2706;
 buffer[578] = 16'h616E;
 buffer[579] = 16'h656D;
 buffer[580] = 16'h003F;
 buffer[581] = 16'hFEB8;
 buffer[582] = 16'h700C;
 buffer[583] = 16'h0482;
 buffer[584] = 16'h2704;
 buffer[585] = 16'h2C24;
 buffer[586] = 16'h006E;
 buffer[587] = 16'hFEBA;
 buffer[588] = 16'h700C;
 buffer[589] = 16'h0490;
 buffer[590] = 16'h2706;
 buffer[591] = 16'h766F;
 buffer[592] = 16'h7265;
 buffer[593] = 16'h0074;
 buffer[594] = 16'hFEBC;
 buffer[595] = 16'h700C;
 buffer[596] = 16'h049C;
 buffer[597] = 16'h2702;
 buffer[598] = 16'h003B;
 buffer[599] = 16'hFEBE;
 buffer[600] = 16'h700C;
 buffer[601] = 16'h04AA;
 buffer[602] = 16'h2707;
 buffer[603] = 16'h7263;
 buffer[604] = 16'h6165;
 buffer[605] = 16'h6574;
 buffer[606] = 16'hFEC0;
 buffer[607] = 16'h700C;
 buffer[608] = 16'h04B4;
 buffer[609] = 16'h3F04;
 buffer[610] = 16'h7564;
 buffer[611] = 16'h0070;
 buffer[612] = 16'h6081;
 buffer[613] = 16'h2267;
 buffer[614] = 16'h708D;
 buffer[615] = 16'h700C;
 buffer[616] = 16'h04C2;
 buffer[617] = 16'h7203;
 buffer[618] = 16'h746F;
 buffer[619] = 16'h6147;
 buffer[620] = 16'h6180;
 buffer[621] = 16'h6B8D;
 buffer[622] = 16'h718C;
 buffer[623] = 16'h04D2;
 buffer[624] = 16'h3205;
 buffer[625] = 16'h7264;
 buffer[626] = 16'h706F;
 buffer[627] = 16'h6103;
 buffer[628] = 16'h710F;
 buffer[629] = 16'h04E0;
 buffer[630] = 16'h3204;
 buffer[631] = 16'h7564;
 buffer[632] = 16'h0070;
 buffer[633] = 16'h6181;
 buffer[634] = 16'h718D;
 buffer[635] = 16'h04EC;
 buffer[636] = 16'h6E06;
 buffer[637] = 16'h6765;
 buffer[638] = 16'h7461;
 buffer[639] = 16'h0065;
 buffer[640] = 16'h7D1C;
 buffer[641] = 16'h04F8;
 buffer[642] = 16'h6407;
 buffer[643] = 16'h656E;
 buffer[644] = 16'h6167;
 buffer[645] = 16'h6574;
 buffer[646] = 16'h6600;
 buffer[647] = 16'h6147;
 buffer[648] = 16'h6600;
 buffer[649] = 16'h8001;
 buffer[650] = 16'h41AB;
 buffer[651] = 16'h6B8D;
 buffer[652] = 16'h720F;
 buffer[653] = 16'h0504;
 buffer[654] = 16'h2D01;
 buffer[655] = 16'h6D10;
 buffer[656] = 16'h720F;
 buffer[657] = 16'h051C;
 buffer[658] = 16'h6103;
 buffer[659] = 16'h7362;
 buffer[660] = 16'h7A1C;
 buffer[661] = 16'h0524;
 buffer[662] = 16'h6D03;
 buffer[663] = 16'h7861;
 buffer[664] = 16'h7B1F;
 buffer[665] = 16'h052C;
 buffer[666] = 16'h6D03;
 buffer[667] = 16'h6E69;
 buffer[668] = 16'h7C1F;
 buffer[669] = 16'h0534;
 buffer[670] = 16'h7706;
 buffer[671] = 16'h7469;
 buffer[672] = 16'h6968;
 buffer[673] = 16'h006E;
 buffer[674] = 16'h6181;
 buffer[675] = 16'h428F;
 buffer[676] = 16'h6147;
 buffer[677] = 16'h428F;
 buffer[678] = 16'h6B8D;
 buffer[679] = 16'h7F0F;
 buffer[680] = 16'h053C;
 buffer[681] = 16'h7506;
 buffer[682] = 16'h2F6D;
 buffer[683] = 16'h6F6D;
 buffer[684] = 16'h0064;
 buffer[685] = 16'h4279;
 buffer[686] = 16'h6F03;
 buffer[687] = 16'h22D6;
 buffer[688] = 16'h6D10;
 buffer[689] = 16'h800F;
 buffer[690] = 16'h6147;
 buffer[691] = 16'h6147;
 buffer[692] = 16'h6081;
 buffer[693] = 16'h41AB;
 buffer[694] = 16'h6147;
 buffer[695] = 16'h6147;
 buffer[696] = 16'h6081;
 buffer[697] = 16'h41AB;
 buffer[698] = 16'h6B8D;
 buffer[699] = 16'h6203;
 buffer[700] = 16'h6081;
 buffer[701] = 16'h6B8D;
 buffer[702] = 16'h6B81;
 buffer[703] = 16'h6180;
 buffer[704] = 16'h6147;
 buffer[705] = 16'h41AB;
 buffer[706] = 16'h6B8D;
 buffer[707] = 16'h6403;
 buffer[708] = 16'h22CA;
 buffer[709] = 16'h6147;
 buffer[710] = 16'h6103;
 buffer[711] = 16'h6310;
 buffer[712] = 16'h6B8D;
 buffer[713] = 16'h02CB;
 buffer[714] = 16'h6103;
 buffer[715] = 16'h6B8D;
 buffer[716] = 16'h6B81;
 buffer[717] = 16'h22D2;
 buffer[718] = 16'h6B8D;
 buffer[719] = 16'h6A00;
 buffer[720] = 16'h6147;
 buffer[721] = 16'h02B3;
 buffer[722] = 16'h6B8D;
 buffer[723] = 16'h6103;
 buffer[724] = 16'h6103;
 buffer[725] = 16'h718C;
 buffer[726] = 16'h6103;
 buffer[727] = 16'h4273;
 buffer[728] = 16'h8000;
 buffer[729] = 16'h6600;
 buffer[730] = 16'h708D;
 buffer[731] = 16'h0552;
 buffer[732] = 16'h6D05;
 buffer[733] = 16'h6D2F;
 buffer[734] = 16'h646F;
 buffer[735] = 16'h6081;
 buffer[736] = 16'h6810;
 buffer[737] = 16'h6081;
 buffer[738] = 16'h6147;
 buffer[739] = 16'h22E8;
 buffer[740] = 16'h6D10;
 buffer[741] = 16'h6147;
 buffer[742] = 16'h4286;
 buffer[743] = 16'h6B8D;
 buffer[744] = 16'h6147;
 buffer[745] = 16'h6081;
 buffer[746] = 16'h6810;
 buffer[747] = 16'h22EE;
 buffer[748] = 16'h6B81;
 buffer[749] = 16'h6203;
 buffer[750] = 16'h6B8D;
 buffer[751] = 16'h42AD;
 buffer[752] = 16'h6B8D;
 buffer[753] = 16'h22F5;
 buffer[754] = 16'h6180;
 buffer[755] = 16'h6D10;
 buffer[756] = 16'h718C;
 buffer[757] = 16'h700C;
 buffer[758] = 16'h05B8;
 buffer[759] = 16'h2F04;
 buffer[760] = 16'h6F6D;
 buffer[761] = 16'h0064;
 buffer[762] = 16'h6181;
 buffer[763] = 16'h6810;
 buffer[764] = 16'h6180;
 buffer[765] = 16'h02DF;
 buffer[766] = 16'h05EE;
 buffer[767] = 16'h6D03;
 buffer[768] = 16'h646F;
 buffer[769] = 16'h42FA;
 buffer[770] = 16'h710F;
 buffer[771] = 16'h05FE;
 buffer[772] = 16'h2F01;
 buffer[773] = 16'h42FA;
 buffer[774] = 16'h700F;
 buffer[775] = 16'h0608;
 buffer[776] = 16'h7503;
 buffer[777] = 16'h2A6D;
 buffer[778] = 16'h8000;
 buffer[779] = 16'h6180;
 buffer[780] = 16'h800F;
 buffer[781] = 16'h6147;
 buffer[782] = 16'h6081;
 buffer[783] = 16'h41AB;
 buffer[784] = 16'h6147;
 buffer[785] = 16'h6147;
 buffer[786] = 16'h6081;
 buffer[787] = 16'h41AB;
 buffer[788] = 16'h6B8D;
 buffer[789] = 16'h6203;
 buffer[790] = 16'h6B8D;
 buffer[791] = 16'h231D;
 buffer[792] = 16'h6147;
 buffer[793] = 16'h6181;
 buffer[794] = 16'h41AB;
 buffer[795] = 16'h6B8D;
 buffer[796] = 16'h6203;
 buffer[797] = 16'h6B81;
 buffer[798] = 16'h2323;
 buffer[799] = 16'h6B8D;
 buffer[800] = 16'h6A00;
 buffer[801] = 16'h6147;
 buffer[802] = 16'h030E;
 buffer[803] = 16'h6B8D;
 buffer[804] = 16'h6103;
 buffer[805] = 16'h426B;
 buffer[806] = 16'h710F;
 buffer[807] = 16'h0610;
 buffer[808] = 16'h2A01;
 buffer[809] = 16'h430A;
 buffer[810] = 16'h710F;
 buffer[811] = 16'h0650;
 buffer[812] = 16'h6D02;
 buffer[813] = 16'h002A;
 buffer[814] = 16'h4279;
 buffer[815] = 16'h6503;
 buffer[816] = 16'h6810;
 buffer[817] = 16'h6147;
 buffer[818] = 16'h6A10;
 buffer[819] = 16'h6180;
 buffer[820] = 16'h6A10;
 buffer[821] = 16'h430A;
 buffer[822] = 16'h6B8D;
 buffer[823] = 16'h2339;
 buffer[824] = 16'h0286;
 buffer[825] = 16'h700C;
 buffer[826] = 16'h0658;
 buffer[827] = 16'h2A05;
 buffer[828] = 16'h6D2F;
 buffer[829] = 16'h646F;
 buffer[830] = 16'h6147;
 buffer[831] = 16'h432E;
 buffer[832] = 16'h6B8D;
 buffer[833] = 16'h02DF;
 buffer[834] = 16'h0676;
 buffer[835] = 16'h2A02;
 buffer[836] = 16'h002F;
 buffer[837] = 16'h433E;
 buffer[838] = 16'h700F;
 buffer[839] = 16'h0686;
 buffer[840] = 16'h6305;
 buffer[841] = 16'h6C65;
 buffer[842] = 16'h2B6C;
 buffer[843] = 16'h8002;
 buffer[844] = 16'h720F;
 buffer[845] = 16'h0690;
 buffer[846] = 16'h6305;
 buffer[847] = 16'h6C65;
 buffer[848] = 16'h2D6C;
 buffer[849] = 16'h8002;
 buffer[850] = 16'h028F;
 buffer[851] = 16'h069C;
 buffer[852] = 16'h6305;
 buffer[853] = 16'h6C65;
 buffer[854] = 16'h736C;
 buffer[855] = 16'h8001;
 buffer[856] = 16'h7D0F;
 buffer[857] = 16'h06A8;
 buffer[858] = 16'h6202;
 buffer[859] = 16'h006C;
 buffer[860] = 16'h8020;
 buffer[861] = 16'h700C;
 buffer[862] = 16'h06B4;
 buffer[863] = 16'h3E05;
 buffer[864] = 16'h6863;
 buffer[865] = 16'h7261;
 buffer[866] = 16'h807F;
 buffer[867] = 16'h6303;
 buffer[868] = 16'h6081;
 buffer[869] = 16'h807F;
 buffer[870] = 16'h435C;
 buffer[871] = 16'h42A2;
 buffer[872] = 16'h236B;
 buffer[873] = 16'h6103;
 buffer[874] = 16'h805F;
 buffer[875] = 16'h700C;
 buffer[876] = 16'h700C;
 buffer[877] = 16'h06BE;
 buffer[878] = 16'h2B02;
 buffer[879] = 16'h0021;
 buffer[880] = 16'h414F;
 buffer[881] = 16'h6C00;
 buffer[882] = 16'h6203;
 buffer[883] = 16'h6180;
 buffer[884] = 16'h6023;
 buffer[885] = 16'h710F;
 buffer[886] = 16'h06DC;
 buffer[887] = 16'h3202;
 buffer[888] = 16'h0021;
 buffer[889] = 16'h6180;
 buffer[890] = 16'h6181;
 buffer[891] = 16'h6023;
 buffer[892] = 16'h6103;
 buffer[893] = 16'h434B;
 buffer[894] = 16'h6023;
 buffer[895] = 16'h710F;
 buffer[896] = 16'h06EE;
 buffer[897] = 16'h3202;
 buffer[898] = 16'h0040;
 buffer[899] = 16'h6081;
 buffer[900] = 16'h434B;
 buffer[901] = 16'h6C00;
 buffer[902] = 16'h6180;
 buffer[903] = 16'h7C0C;
 buffer[904] = 16'h0702;
 buffer[905] = 16'h6305;
 buffer[906] = 16'h756F;
 buffer[907] = 16'h746E;
 buffer[908] = 16'h6081;
 buffer[909] = 16'h6310;
 buffer[910] = 16'h6180;
 buffer[911] = 16'h017E;
 buffer[912] = 16'h0712;
 buffer[913] = 16'h6804;
 buffer[914] = 16'h7265;
 buffer[915] = 16'h0065;
 buffer[916] = 16'hFEAC;
 buffer[917] = 16'h7C0C;
 buffer[918] = 16'h0722;
 buffer[919] = 16'h6107;
 buffer[920] = 16'h696C;
 buffer[921] = 16'h6E67;
 buffer[922] = 16'h6465;
 buffer[923] = 16'h6081;
 buffer[924] = 16'h8000;
 buffer[925] = 16'h8002;
 buffer[926] = 16'h42AD;
 buffer[927] = 16'h6103;
 buffer[928] = 16'h6081;
 buffer[929] = 16'h23A5;
 buffer[930] = 16'h8002;
 buffer[931] = 16'h6180;
 buffer[932] = 16'h428F;
 buffer[933] = 16'h720F;
 buffer[934] = 16'h072E;
 buffer[935] = 16'h6105;
 buffer[936] = 16'h696C;
 buffer[937] = 16'h6E67;
 buffer[938] = 16'h4394;
 buffer[939] = 16'h439B;
 buffer[940] = 16'hFEAC;
 buffer[941] = 16'h6023;
 buffer[942] = 16'h710F;
 buffer[943] = 16'h074E;
 buffer[944] = 16'h7003;
 buffer[945] = 16'h6461;
 buffer[946] = 16'h4394;
 buffer[947] = 16'h8050;
 buffer[948] = 16'h6203;
 buffer[949] = 16'h039B;
 buffer[950] = 16'h0760;
 buffer[951] = 16'h4008;
 buffer[952] = 16'h7865;
 buffer[953] = 16'h6365;
 buffer[954] = 16'h7475;
 buffer[955] = 16'h0065;
 buffer[956] = 16'h6C00;
 buffer[957] = 16'h4264;
 buffer[958] = 16'h23C0;
 buffer[959] = 16'h0172;
 buffer[960] = 16'h700C;
 buffer[961] = 16'h076E;
 buffer[962] = 16'h6604;
 buffer[963] = 16'h6C69;
 buffer[964] = 16'h006C;
 buffer[965] = 16'h6180;
 buffer[966] = 16'h6147;
 buffer[967] = 16'h6180;
 buffer[968] = 16'h03CC;
 buffer[969] = 16'h4279;
 buffer[970] = 16'h418D;
 buffer[971] = 16'h6310;
 buffer[972] = 16'h6B81;
 buffer[973] = 16'h23D2;
 buffer[974] = 16'h6B8D;
 buffer[975] = 16'h6A00;
 buffer[976] = 16'h6147;
 buffer[977] = 16'h03C9;
 buffer[978] = 16'h6B8D;
 buffer[979] = 16'h6103;
 buffer[980] = 16'h0273;
 buffer[981] = 16'h0784;
 buffer[982] = 16'h6505;
 buffer[983] = 16'h6172;
 buffer[984] = 16'h6573;
 buffer[985] = 16'h8000;
 buffer[986] = 16'h03C5;
 buffer[987] = 16'h07AC;
 buffer[988] = 16'h6405;
 buffer[989] = 16'h6769;
 buffer[990] = 16'h7469;
 buffer[991] = 16'h8009;
 buffer[992] = 16'h6181;
 buffer[993] = 16'h6803;
 buffer[994] = 16'h8007;
 buffer[995] = 16'h6303;
 buffer[996] = 16'h6203;
 buffer[997] = 16'h8030;
 buffer[998] = 16'h720F;
 buffer[999] = 16'h07B8;
 buffer[1000] = 16'h6507;
 buffer[1001] = 16'h7478;
 buffer[1002] = 16'h6172;
 buffer[1003] = 16'h7463;
 buffer[1004] = 16'h8000;
 buffer[1005] = 16'h6180;
 buffer[1006] = 16'h42AD;
 buffer[1007] = 16'h6180;
 buffer[1008] = 16'h03DF;
 buffer[1009] = 16'h07D0;
 buffer[1010] = 16'h3C02;
 buffer[1011] = 16'h0023;
 buffer[1012] = 16'h43B2;
 buffer[1013] = 16'hFE8E;
 buffer[1014] = 16'h6023;
 buffer[1015] = 16'h710F;
 buffer[1016] = 16'h07E4;
 buffer[1017] = 16'h6804;
 buffer[1018] = 16'h6C6F;
 buffer[1019] = 16'h0064;
 buffer[1020] = 16'hFE8E;
 buffer[1021] = 16'h6C00;
 buffer[1022] = 16'h6A00;
 buffer[1023] = 16'h6081;
 buffer[1024] = 16'hFE8E;
 buffer[1025] = 16'h6023;
 buffer[1026] = 16'h6103;
 buffer[1027] = 16'h018D;
 buffer[1028] = 16'h07F2;
 buffer[1029] = 16'h2301;
 buffer[1030] = 16'hFE80;
 buffer[1031] = 16'h6C00;
 buffer[1032] = 16'h43EC;
 buffer[1033] = 16'h03FC;
 buffer[1034] = 16'h080A;
 buffer[1035] = 16'h2302;
 buffer[1036] = 16'h0073;
 buffer[1037] = 16'h4406;
 buffer[1038] = 16'h6081;
 buffer[1039] = 16'h2411;
 buffer[1040] = 16'h040D;
 buffer[1041] = 16'h700C;
 buffer[1042] = 16'h0816;
 buffer[1043] = 16'h7304;
 buffer[1044] = 16'h6769;
 buffer[1045] = 16'h006E;
 buffer[1046] = 16'h6810;
 buffer[1047] = 16'h241A;
 buffer[1048] = 16'h802D;
 buffer[1049] = 16'h03FC;
 buffer[1050] = 16'h700C;
 buffer[1051] = 16'h0826;
 buffer[1052] = 16'h2302;
 buffer[1053] = 16'h003E;
 buffer[1054] = 16'h6103;
 buffer[1055] = 16'hFE8E;
 buffer[1056] = 16'h6C00;
 buffer[1057] = 16'h43B2;
 buffer[1058] = 16'h6181;
 buffer[1059] = 16'h028F;
 buffer[1060] = 16'h0838;
 buffer[1061] = 16'h7303;
 buffer[1062] = 16'h7274;
 buffer[1063] = 16'h6081;
 buffer[1064] = 16'h6147;
 buffer[1065] = 16'h6A10;
 buffer[1066] = 16'h43F4;
 buffer[1067] = 16'h440D;
 buffer[1068] = 16'h6B8D;
 buffer[1069] = 16'h4416;
 buffer[1070] = 16'h041E;
 buffer[1071] = 16'h084A;
 buffer[1072] = 16'h6803;
 buffer[1073] = 16'h7865;
 buffer[1074] = 16'h8010;
 buffer[1075] = 16'hFE80;
 buffer[1076] = 16'h6023;
 buffer[1077] = 16'h710F;
 buffer[1078] = 16'h0860;
 buffer[1079] = 16'h6407;
 buffer[1080] = 16'h6365;
 buffer[1081] = 16'h6D69;
 buffer[1082] = 16'h6C61;
 buffer[1083] = 16'h800A;
 buffer[1084] = 16'hFE80;
 buffer[1085] = 16'h6023;
 buffer[1086] = 16'h710F;
 buffer[1087] = 16'h086E;
 buffer[1088] = 16'h6406;
 buffer[1089] = 16'h6769;
 buffer[1090] = 16'h7469;
 buffer[1091] = 16'h003F;
 buffer[1092] = 16'h6147;
 buffer[1093] = 16'h8030;
 buffer[1094] = 16'h428F;
 buffer[1095] = 16'h8009;
 buffer[1096] = 16'h6181;
 buffer[1097] = 16'h6803;
 buffer[1098] = 16'h2457;
 buffer[1099] = 16'h6081;
 buffer[1100] = 16'h8020;
 buffer[1101] = 16'h6613;
 buffer[1102] = 16'h2451;
 buffer[1103] = 16'h8020;
 buffer[1104] = 16'h428F;
 buffer[1105] = 16'h8007;
 buffer[1106] = 16'h428F;
 buffer[1107] = 16'h6081;
 buffer[1108] = 16'h800A;
 buffer[1109] = 16'h6803;
 buffer[1110] = 16'h6403;
 buffer[1111] = 16'h6081;
 buffer[1112] = 16'h6B8D;
 buffer[1113] = 16'h7F0F;
 buffer[1114] = 16'h0880;
 buffer[1115] = 16'h6E07;
 buffer[1116] = 16'h6D75;
 buffer[1117] = 16'h6562;
 buffer[1118] = 16'h3F72;
 buffer[1119] = 16'hFE80;
 buffer[1120] = 16'h6C00;
 buffer[1121] = 16'h6147;
 buffer[1122] = 16'h8000;
 buffer[1123] = 16'h6181;
 buffer[1124] = 16'h438C;
 buffer[1125] = 16'h6181;
 buffer[1126] = 16'h417E;
 buffer[1127] = 16'h8024;
 buffer[1128] = 16'h6703;
 buffer[1129] = 16'h246F;
 buffer[1130] = 16'h4432;
 buffer[1131] = 16'h6180;
 buffer[1132] = 16'h6310;
 buffer[1133] = 16'h6180;
 buffer[1134] = 16'h6A00;
 buffer[1135] = 16'h6181;
 buffer[1136] = 16'h417E;
 buffer[1137] = 16'h802D;
 buffer[1138] = 16'h6703;
 buffer[1139] = 16'h6147;
 buffer[1140] = 16'h6180;
 buffer[1141] = 16'h6B81;
 buffer[1142] = 16'h428F;
 buffer[1143] = 16'h6180;
 buffer[1144] = 16'h6B81;
 buffer[1145] = 16'h6203;
 buffer[1146] = 16'h4264;
 buffer[1147] = 16'h24A0;
 buffer[1148] = 16'h6A00;
 buffer[1149] = 16'h6147;
 buffer[1150] = 16'h6081;
 buffer[1151] = 16'h6147;
 buffer[1152] = 16'h417E;
 buffer[1153] = 16'hFE80;
 buffer[1154] = 16'h6C00;
 buffer[1155] = 16'h4444;
 buffer[1156] = 16'h249A;
 buffer[1157] = 16'h6180;
 buffer[1158] = 16'hFE80;
 buffer[1159] = 16'h6C00;
 buffer[1160] = 16'h4329;
 buffer[1161] = 16'h6203;
 buffer[1162] = 16'h6B8D;
 buffer[1163] = 16'h6310;
 buffer[1164] = 16'h6B81;
 buffer[1165] = 16'h2492;
 buffer[1166] = 16'h6B8D;
 buffer[1167] = 16'h6A00;
 buffer[1168] = 16'h6147;
 buffer[1169] = 16'h047E;
 buffer[1170] = 16'h6B8D;
 buffer[1171] = 16'h6103;
 buffer[1172] = 16'h6B81;
 buffer[1173] = 16'h6003;
 buffer[1174] = 16'h2498;
 buffer[1175] = 16'h6D10;
 buffer[1176] = 16'h6180;
 buffer[1177] = 16'h049F;
 buffer[1178] = 16'h6B8D;
 buffer[1179] = 16'h6B8D;
 buffer[1180] = 16'h4273;
 buffer[1181] = 16'h4273;
 buffer[1182] = 16'h8000;
 buffer[1183] = 16'h6081;
 buffer[1184] = 16'h6B8D;
 buffer[1185] = 16'h4273;
 buffer[1186] = 16'h6B8D;
 buffer[1187] = 16'hFE80;
 buffer[1188] = 16'h6023;
 buffer[1189] = 16'h710F;
 buffer[1190] = 16'h08B6;
 buffer[1191] = 16'h3F03;
 buffer[1192] = 16'h7872;
 buffer[1193] = 16'h8FFE;
 buffer[1194] = 16'h6600;
 buffer[1195] = 16'h6C00;
 buffer[1196] = 16'h8001;
 buffer[1197] = 16'h6303;
 buffer[1198] = 16'h711C;
 buffer[1199] = 16'h094E;
 buffer[1200] = 16'h7403;
 buffer[1201] = 16'h2178;
 buffer[1202] = 16'h8FFE;
 buffer[1203] = 16'h6600;
 buffer[1204] = 16'h6C00;
 buffer[1205] = 16'h8002;
 buffer[1206] = 16'h6303;
 buffer[1207] = 16'h6010;
 buffer[1208] = 16'h24B2;
 buffer[1209] = 16'h6081;
 buffer[1210] = 16'h8FFF;
 buffer[1211] = 16'h6600;
 buffer[1212] = 16'h6023;
 buffer[1213] = 16'h6103;
 buffer[1214] = 16'h80DF;
 buffer[1215] = 16'h6600;
 buffer[1216] = 16'h6023;
 buffer[1217] = 16'h710F;
 buffer[1218] = 16'h0960;
 buffer[1219] = 16'h3F04;
 buffer[1220] = 16'h656B;
 buffer[1221] = 16'h0079;
 buffer[1222] = 16'hFEB0;
 buffer[1223] = 16'h03BC;
 buffer[1224] = 16'h0986;
 buffer[1225] = 16'h6504;
 buffer[1226] = 16'h696D;
 buffer[1227] = 16'h0074;
 buffer[1228] = 16'hFEB2;
 buffer[1229] = 16'h03BC;
 buffer[1230] = 16'h0992;
 buffer[1231] = 16'h6B03;
 buffer[1232] = 16'h7965;
 buffer[1233] = 16'h44C6;
 buffer[1234] = 16'h24D1;
 buffer[1235] = 16'h8FFF;
 buffer[1236] = 16'h6600;
 buffer[1237] = 16'h7C0C;
 buffer[1238] = 16'h099E;
 buffer[1239] = 16'h6E04;
 buffer[1240] = 16'h6675;
 buffer[1241] = 16'h003F;
 buffer[1242] = 16'h44C6;
 buffer[1243] = 16'h6081;
 buffer[1244] = 16'h24E1;
 buffer[1245] = 16'h6103;
 buffer[1246] = 16'h44D1;
 buffer[1247] = 16'h800D;
 buffer[1248] = 16'h770F;
 buffer[1249] = 16'h700C;
 buffer[1250] = 16'h09AE;
 buffer[1251] = 16'h7406;
 buffer[1252] = 16'h6D69;
 buffer[1253] = 16'h7265;
 buffer[1254] = 16'h0040;
 buffer[1255] = 16'h8FFB;
 buffer[1256] = 16'h6600;
 buffer[1257] = 16'h7C0C;
 buffer[1258] = 16'h09C6;
 buffer[1259] = 16'h6C04;
 buffer[1260] = 16'h6465;
 buffer[1261] = 16'h0040;
 buffer[1262] = 16'h8FFD;
 buffer[1263] = 16'h6600;
 buffer[1264] = 16'h7C0C;
 buffer[1265] = 16'h09D6;
 buffer[1266] = 16'h6C04;
 buffer[1267] = 16'h6465;
 buffer[1268] = 16'h0021;
 buffer[1269] = 16'h8FFD;
 buffer[1270] = 16'h6600;
 buffer[1271] = 16'h6023;
 buffer[1272] = 16'h710F;
 buffer[1273] = 16'h09E4;
 buffer[1274] = 16'h6208;
 buffer[1275] = 16'h7475;
 buffer[1276] = 16'h6F74;
 buffer[1277] = 16'h736E;
 buffer[1278] = 16'h0040;
 buffer[1279] = 16'h8FFC;
 buffer[1280] = 16'h6600;
 buffer[1281] = 16'h7C0C;
 buffer[1282] = 16'h09F4;
 buffer[1283] = 16'h7305;
 buffer[1284] = 16'h6170;
 buffer[1285] = 16'h6563;
 buffer[1286] = 16'h435C;
 buffer[1287] = 16'h04CC;
 buffer[1288] = 16'h0A06;
 buffer[1289] = 16'h7306;
 buffer[1290] = 16'h6170;
 buffer[1291] = 16'h6563;
 buffer[1292] = 16'h0073;
 buffer[1293] = 16'h8000;
 buffer[1294] = 16'h6B13;
 buffer[1295] = 16'h6147;
 buffer[1296] = 16'h0512;
 buffer[1297] = 16'h4506;
 buffer[1298] = 16'h6B81;
 buffer[1299] = 16'h2518;
 buffer[1300] = 16'h6B8D;
 buffer[1301] = 16'h6A00;
 buffer[1302] = 16'h6147;
 buffer[1303] = 16'h0511;
 buffer[1304] = 16'h6B8D;
 buffer[1305] = 16'h710F;
 buffer[1306] = 16'h0A12;
 buffer[1307] = 16'h7404;
 buffer[1308] = 16'h7079;
 buffer[1309] = 16'h0065;
 buffer[1310] = 16'h6147;
 buffer[1311] = 16'h0522;
 buffer[1312] = 16'h438C;
 buffer[1313] = 16'h44CC;
 buffer[1314] = 16'h6B81;
 buffer[1315] = 16'h2528;
 buffer[1316] = 16'h6B8D;
 buffer[1317] = 16'h6A00;
 buffer[1318] = 16'h6147;
 buffer[1319] = 16'h0520;
 buffer[1320] = 16'h6B8D;
 buffer[1321] = 16'h6103;
 buffer[1322] = 16'h710F;
 buffer[1323] = 16'h0A36;
 buffer[1324] = 16'h6302;
 buffer[1325] = 16'h0072;
 buffer[1326] = 16'h800D;
 buffer[1327] = 16'h44CC;
 buffer[1328] = 16'h800A;
 buffer[1329] = 16'h04CC;
 buffer[1330] = 16'h0A58;
 buffer[1331] = 16'h6443;
 buffer[1332] = 16'h246F;
 buffer[1333] = 16'h6B8D;
 buffer[1334] = 16'h6B81;
 buffer[1335] = 16'h6B8D;
 buffer[1336] = 16'h438C;
 buffer[1337] = 16'h6203;
 buffer[1338] = 16'h439B;
 buffer[1339] = 16'h6147;
 buffer[1340] = 16'h6180;
 buffer[1341] = 16'h6147;
 buffer[1342] = 16'h700C;
 buffer[1343] = 16'h0A66;
 buffer[1344] = 16'h2443;
 buffer[1345] = 16'h7C22;
 buffer[1346] = 16'h4535;
 buffer[1347] = 16'h700C;
 buffer[1348] = 16'h0A80;
 buffer[1349] = 16'h2E02;
 buffer[1350] = 16'h0024;
 buffer[1351] = 16'h438C;
 buffer[1352] = 16'h051E;
 buffer[1353] = 16'h0A8A;
 buffer[1354] = 16'h2E43;
 buffer[1355] = 16'h7C22;
 buffer[1356] = 16'h4535;
 buffer[1357] = 16'h0547;
 buffer[1358] = 16'h0A94;
 buffer[1359] = 16'h2E02;
 buffer[1360] = 16'h0072;
 buffer[1361] = 16'h6147;
 buffer[1362] = 16'h4427;
 buffer[1363] = 16'h6B8D;
 buffer[1364] = 16'h6181;
 buffer[1365] = 16'h428F;
 buffer[1366] = 16'h450D;
 buffer[1367] = 16'h051E;
 buffer[1368] = 16'h0A9E;
 buffer[1369] = 16'h7503;
 buffer[1370] = 16'h722E;
 buffer[1371] = 16'h6147;
 buffer[1372] = 16'h43F4;
 buffer[1373] = 16'h440D;
 buffer[1374] = 16'h441E;
 buffer[1375] = 16'h6B8D;
 buffer[1376] = 16'h6181;
 buffer[1377] = 16'h428F;
 buffer[1378] = 16'h450D;
 buffer[1379] = 16'h051E;
 buffer[1380] = 16'h0AB2;
 buffer[1381] = 16'h7502;
 buffer[1382] = 16'h002E;
 buffer[1383] = 16'h43F4;
 buffer[1384] = 16'h440D;
 buffer[1385] = 16'h441E;
 buffer[1386] = 16'h4506;
 buffer[1387] = 16'h051E;
 buffer[1388] = 16'h0ACA;
 buffer[1389] = 16'h2E01;
 buffer[1390] = 16'hFE80;
 buffer[1391] = 16'h6C00;
 buffer[1392] = 16'h800A;
 buffer[1393] = 16'h6503;
 buffer[1394] = 16'h2574;
 buffer[1395] = 16'h0567;
 buffer[1396] = 16'h4427;
 buffer[1397] = 16'h4506;
 buffer[1398] = 16'h051E;
 buffer[1399] = 16'h0ADA;
 buffer[1400] = 16'h2E02;
 buffer[1401] = 16'h0023;
 buffer[1402] = 16'hFE80;
 buffer[1403] = 16'h6C00;
 buffer[1404] = 16'h6180;
 buffer[1405] = 16'h443B;
 buffer[1406] = 16'h456E;
 buffer[1407] = 16'hFE80;
 buffer[1408] = 16'h6023;
 buffer[1409] = 16'h710F;
 buffer[1410] = 16'h0AF0;
 buffer[1411] = 16'h7503;
 buffer[1412] = 16'h232E;
 buffer[1413] = 16'hFE80;
 buffer[1414] = 16'h6C00;
 buffer[1415] = 16'h6180;
 buffer[1416] = 16'h443B;
 buffer[1417] = 16'h43F4;
 buffer[1418] = 16'h440D;
 buffer[1419] = 16'h441E;
 buffer[1420] = 16'h4506;
 buffer[1421] = 16'h451E;
 buffer[1422] = 16'hFE80;
 buffer[1423] = 16'h6023;
 buffer[1424] = 16'h710F;
 buffer[1425] = 16'h0B06;
 buffer[1426] = 16'h7504;
 buffer[1427] = 16'h722E;
 buffer[1428] = 16'h0023;
 buffer[1429] = 16'hFE80;
 buffer[1430] = 16'h6C00;
 buffer[1431] = 16'h426B;
 buffer[1432] = 16'h426B;
 buffer[1433] = 16'h443B;
 buffer[1434] = 16'h6147;
 buffer[1435] = 16'h43F4;
 buffer[1436] = 16'h440D;
 buffer[1437] = 16'h441E;
 buffer[1438] = 16'h6B8D;
 buffer[1439] = 16'h6181;
 buffer[1440] = 16'h428F;
 buffer[1441] = 16'h450D;
 buffer[1442] = 16'h451E;
 buffer[1443] = 16'hFE80;
 buffer[1444] = 16'h6023;
 buffer[1445] = 16'h710F;
 buffer[1446] = 16'h0B24;
 buffer[1447] = 16'h2E03;
 buffer[1448] = 16'h2372;
 buffer[1449] = 16'hFE80;
 buffer[1450] = 16'h6C00;
 buffer[1451] = 16'h426B;
 buffer[1452] = 16'h426B;
 buffer[1453] = 16'h443B;
 buffer[1454] = 16'h6147;
 buffer[1455] = 16'h4427;
 buffer[1456] = 16'h6B8D;
 buffer[1457] = 16'h6181;
 buffer[1458] = 16'h428F;
 buffer[1459] = 16'h450D;
 buffer[1460] = 16'h451E;
 buffer[1461] = 16'hFE80;
 buffer[1462] = 16'h6023;
 buffer[1463] = 16'h710F;
 buffer[1464] = 16'h0B4E;
 buffer[1465] = 16'h6305;
 buffer[1466] = 16'h6F6D;
 buffer[1467] = 16'h6576;
 buffer[1468] = 16'h6147;
 buffer[1469] = 16'h05C6;
 buffer[1470] = 16'h6147;
 buffer[1471] = 16'h6081;
 buffer[1472] = 16'h417E;
 buffer[1473] = 16'h6B81;
 buffer[1474] = 16'h418D;
 buffer[1475] = 16'h6310;
 buffer[1476] = 16'h6B8D;
 buffer[1477] = 16'h6310;
 buffer[1478] = 16'h6B81;
 buffer[1479] = 16'h25CC;
 buffer[1480] = 16'h6B8D;
 buffer[1481] = 16'h6A00;
 buffer[1482] = 16'h6147;
 buffer[1483] = 16'h05BE;
 buffer[1484] = 16'h6B8D;
 buffer[1485] = 16'h6103;
 buffer[1486] = 16'h0273;
 buffer[1487] = 16'h0B72;
 buffer[1488] = 16'h7005;
 buffer[1489] = 16'h6361;
 buffer[1490] = 16'h246B;
 buffer[1491] = 16'h6081;
 buffer[1492] = 16'h6147;
 buffer[1493] = 16'h4279;
 buffer[1494] = 16'h6023;
 buffer[1495] = 16'h6103;
 buffer[1496] = 16'h6310;
 buffer[1497] = 16'h6180;
 buffer[1498] = 16'h45BC;
 buffer[1499] = 16'h6B8D;
 buffer[1500] = 16'h700C;
 buffer[1501] = 16'h0BA0;
 buffer[1502] = 16'h3F01;
 buffer[1503] = 16'h6C00;
 buffer[1504] = 16'h056E;
 buffer[1505] = 16'h0BBC;
 buffer[1506] = 16'h3205;
 buffer[1507] = 16'h766F;
 buffer[1508] = 16'h7265;
 buffer[1509] = 16'h6147;
 buffer[1510] = 16'h6147;
 buffer[1511] = 16'h4279;
 buffer[1512] = 16'h6B8D;
 buffer[1513] = 16'h6B8D;
 buffer[1514] = 16'h426B;
 buffer[1515] = 16'h6147;
 buffer[1516] = 16'h426B;
 buffer[1517] = 16'h6B8D;
 buffer[1518] = 16'h700C;
 buffer[1519] = 16'h0BC4;
 buffer[1520] = 16'h3205;
 buffer[1521] = 16'h7773;
 buffer[1522] = 16'h7061;
 buffer[1523] = 16'h426B;
 buffer[1524] = 16'h6147;
 buffer[1525] = 16'h426B;
 buffer[1526] = 16'h6B8D;
 buffer[1527] = 16'h700C;
 buffer[1528] = 16'h0BE0;
 buffer[1529] = 16'h3204;
 buffer[1530] = 16'h696E;
 buffer[1531] = 16'h0070;
 buffer[1532] = 16'h426B;
 buffer[1533] = 16'h6103;
 buffer[1534] = 16'h426B;
 buffer[1535] = 16'h710F;
 buffer[1536] = 16'h0BF2;
 buffer[1537] = 16'h3204;
 buffer[1538] = 16'h6F72;
 buffer[1539] = 16'h0074;
 buffer[1540] = 16'h6180;
 buffer[1541] = 16'h6147;
 buffer[1542] = 16'h6147;
 buffer[1543] = 16'h45F3;
 buffer[1544] = 16'h6B8D;
 buffer[1545] = 16'h6B8D;
 buffer[1546] = 16'h6180;
 buffer[1547] = 16'h05F3;
 buffer[1548] = 16'h0C02;
 buffer[1549] = 16'h6402;
 buffer[1550] = 16'h003D;
 buffer[1551] = 16'h6147;
 buffer[1552] = 16'h426B;
 buffer[1553] = 16'h6503;
 buffer[1554] = 16'h6180;
 buffer[1555] = 16'h6B8D;
 buffer[1556] = 16'h6503;
 buffer[1557] = 16'h6403;
 buffer[1558] = 16'h701C;
 buffer[1559] = 16'h0C1A;
 buffer[1560] = 16'h6403;
 buffer[1561] = 16'h3E3C;
 buffer[1562] = 16'h460F;
 buffer[1563] = 16'h760C;
 buffer[1564] = 16'h0C30;
 buffer[1565] = 16'h6402;
 buffer[1566] = 16'h002B;
 buffer[1567] = 16'h426B;
 buffer[1568] = 16'h6203;
 buffer[1569] = 16'h6147;
 buffer[1570] = 16'h6181;
 buffer[1571] = 16'h6203;
 buffer[1572] = 16'h6081;
 buffer[1573] = 16'h426B;
 buffer[1574] = 16'h6F03;
 buffer[1575] = 16'h262B;
 buffer[1576] = 16'h6B8D;
 buffer[1577] = 16'h6310;
 buffer[1578] = 16'h062C;
 buffer[1579] = 16'h6B8D;
 buffer[1580] = 16'h700C;
 buffer[1581] = 16'h0C3A;
 buffer[1582] = 16'h6402;
 buffer[1583] = 16'h002D;
 buffer[1584] = 16'h4286;
 buffer[1585] = 16'h061F;
 buffer[1586] = 16'h0C5C;
 buffer[1587] = 16'h7303;
 buffer[1588] = 16'h643E;
 buffer[1589] = 16'h6081;
 buffer[1590] = 16'h781C;
 buffer[1591] = 16'h0C66;
 buffer[1592] = 16'h6403;
 buffer[1593] = 16'h2B31;
 buffer[1594] = 16'h8001;
 buffer[1595] = 16'h4635;
 buffer[1596] = 16'h061F;
 buffer[1597] = 16'h0C70;
 buffer[1598] = 16'h6404;
 buffer[1599] = 16'h6F78;
 buffer[1600] = 16'h0072;
 buffer[1601] = 16'h426B;
 buffer[1602] = 16'h6503;
 buffer[1603] = 16'h4155;
 buffer[1604] = 16'h6503;
 buffer[1605] = 16'h718C;
 buffer[1606] = 16'h0C7C;
 buffer[1607] = 16'h6404;
 buffer[1608] = 16'h6E61;
 buffer[1609] = 16'h0064;
 buffer[1610] = 16'h426B;
 buffer[1611] = 16'h6303;
 buffer[1612] = 16'h4155;
 buffer[1613] = 16'h6303;
 buffer[1614] = 16'h718C;
 buffer[1615] = 16'h0C8E;
 buffer[1616] = 16'h6403;
 buffer[1617] = 16'h726F;
 buffer[1618] = 16'h426B;
 buffer[1619] = 16'h6403;
 buffer[1620] = 16'h4155;
 buffer[1621] = 16'h6403;
 buffer[1622] = 16'h718C;
 buffer[1623] = 16'h0CA0;
 buffer[1624] = 16'h6407;
 buffer[1625] = 16'h6E69;
 buffer[1626] = 16'h6576;
 buffer[1627] = 16'h7472;
 buffer[1628] = 16'h6600;
 buffer[1629] = 16'h6180;
 buffer[1630] = 16'h6600;
 buffer[1631] = 16'h718C;
 buffer[1632] = 16'h0CB0;
 buffer[1633] = 16'h6402;
 buffer[1634] = 16'h003C;
 buffer[1635] = 16'h426B;
 buffer[1636] = 16'h4279;
 buffer[1637] = 16'h6703;
 buffer[1638] = 16'h266A;
 buffer[1639] = 16'h4273;
 buffer[1640] = 16'h6F03;
 buffer[1641] = 16'h066C;
 buffer[1642] = 16'h45FC;
 buffer[1643] = 16'h761F;
 buffer[1644] = 16'h0CC2;
 buffer[1645] = 16'h6402;
 buffer[1646] = 16'h003E;
 buffer[1647] = 16'h45F3;
 buffer[1648] = 16'h0663;
 buffer[1649] = 16'h0CDA;
 buffer[1650] = 16'h6403;
 buffer[1651] = 16'h3D30;
 buffer[1652] = 16'h6403;
 buffer[1653] = 16'h701C;
 buffer[1654] = 16'h0CE4;
 buffer[1655] = 16'h6403;
 buffer[1656] = 16'h3C30;
 buffer[1657] = 16'h8000;
 buffer[1658] = 16'h4635;
 buffer[1659] = 16'h0663;
 buffer[1660] = 16'h0CEE;
 buffer[1661] = 16'h6404;
 buffer[1662] = 16'h3C30;
 buffer[1663] = 16'h003E;
 buffer[1664] = 16'h4674;
 buffer[1665] = 16'h760C;
 buffer[1666] = 16'h0CFA;
 buffer[1667] = 16'h6403;
 buffer[1668] = 16'h2A32;
 buffer[1669] = 16'h4279;
 buffer[1670] = 16'h061F;
 buffer[1671] = 16'h0D06;
 buffer[1672] = 16'h6403;
 buffer[1673] = 16'h2F32;
 buffer[1674] = 16'h6081;
 buffer[1675] = 16'h800F;
 buffer[1676] = 16'h6D03;
 buffer[1677] = 16'h6147;
 buffer[1678] = 16'h415D;
 buffer[1679] = 16'h6180;
 buffer[1680] = 16'h415D;
 buffer[1681] = 16'h6B8D;
 buffer[1682] = 16'h6403;
 buffer[1683] = 16'h718C;
 buffer[1684] = 16'h0D10;
 buffer[1685] = 16'h6403;
 buffer[1686] = 16'h2D31;
 buffer[1687] = 16'h8001;
 buffer[1688] = 16'h4635;
 buffer[1689] = 16'h4286;
 buffer[1690] = 16'h061F;
 buffer[1691] = 16'h0D2A;
 buffer[1692] = 16'h2807;
 buffer[1693] = 16'h6170;
 buffer[1694] = 16'h7372;
 buffer[1695] = 16'h2965;
 buffer[1696] = 16'hFE82;
 buffer[1697] = 16'h6023;
 buffer[1698] = 16'h6103;
 buffer[1699] = 16'h6181;
 buffer[1700] = 16'h6147;
 buffer[1701] = 16'h6081;
 buffer[1702] = 16'h26EB;
 buffer[1703] = 16'h6A00;
 buffer[1704] = 16'hFE82;
 buffer[1705] = 16'h6C00;
 buffer[1706] = 16'h435C;
 buffer[1707] = 16'h6703;
 buffer[1708] = 16'h26C7;
 buffer[1709] = 16'h6147;
 buffer[1710] = 16'h438C;
 buffer[1711] = 16'hFE82;
 buffer[1712] = 16'h6C00;
 buffer[1713] = 16'h6180;
 buffer[1714] = 16'h428F;
 buffer[1715] = 16'h6810;
 buffer[1716] = 16'h6600;
 buffer[1717] = 16'h6B81;
 buffer[1718] = 16'h6910;
 buffer[1719] = 16'h6303;
 buffer[1720] = 16'h26C5;
 buffer[1721] = 16'h6B81;
 buffer[1722] = 16'h26BF;
 buffer[1723] = 16'h6B8D;
 buffer[1724] = 16'h6A00;
 buffer[1725] = 16'h6147;
 buffer[1726] = 16'h06AE;
 buffer[1727] = 16'h6B8D;
 buffer[1728] = 16'h6103;
 buffer[1729] = 16'h6B8D;
 buffer[1730] = 16'h6103;
 buffer[1731] = 16'h8000;
 buffer[1732] = 16'h708D;
 buffer[1733] = 16'h6A00;
 buffer[1734] = 16'h6B8D;
 buffer[1735] = 16'h6181;
 buffer[1736] = 16'h6180;
 buffer[1737] = 16'h6147;
 buffer[1738] = 16'h438C;
 buffer[1739] = 16'hFE82;
 buffer[1740] = 16'h6C00;
 buffer[1741] = 16'h6180;
 buffer[1742] = 16'h428F;
 buffer[1743] = 16'hFE82;
 buffer[1744] = 16'h6C00;
 buffer[1745] = 16'h435C;
 buffer[1746] = 16'h6703;
 buffer[1747] = 16'h26D5;
 buffer[1748] = 16'h6810;
 buffer[1749] = 16'h26E1;
 buffer[1750] = 16'h6B81;
 buffer[1751] = 16'h26DC;
 buffer[1752] = 16'h6B8D;
 buffer[1753] = 16'h6A00;
 buffer[1754] = 16'h6147;
 buffer[1755] = 16'h06CA;
 buffer[1756] = 16'h6B8D;
 buffer[1757] = 16'h6103;
 buffer[1758] = 16'h6081;
 buffer[1759] = 16'h6147;
 buffer[1760] = 16'h06E6;
 buffer[1761] = 16'h6B8D;
 buffer[1762] = 16'h6103;
 buffer[1763] = 16'h6081;
 buffer[1764] = 16'h6147;
 buffer[1765] = 16'h6A00;
 buffer[1766] = 16'h6181;
 buffer[1767] = 16'h428F;
 buffer[1768] = 16'h6B8D;
 buffer[1769] = 16'h6B8D;
 buffer[1770] = 16'h028F;
 buffer[1771] = 16'h6181;
 buffer[1772] = 16'h6B8D;
 buffer[1773] = 16'h028F;
 buffer[1774] = 16'h0D38;
 buffer[1775] = 16'h7005;
 buffer[1776] = 16'h7261;
 buffer[1777] = 16'h6573;
 buffer[1778] = 16'h6147;
 buffer[1779] = 16'hFE88;
 buffer[1780] = 16'h6C00;
 buffer[1781] = 16'hFE84;
 buffer[1782] = 16'h6C00;
 buffer[1783] = 16'h6203;
 buffer[1784] = 16'hFE86;
 buffer[1785] = 16'h6C00;
 buffer[1786] = 16'hFE84;
 buffer[1787] = 16'h6C00;
 buffer[1788] = 16'h428F;
 buffer[1789] = 16'h6B8D;
 buffer[1790] = 16'h46A0;
 buffer[1791] = 16'hFE84;
 buffer[1792] = 16'h0370;
 buffer[1793] = 16'h0DDE;
 buffer[1794] = 16'h2E82;
 buffer[1795] = 16'h0028;
 buffer[1796] = 16'h8029;
 buffer[1797] = 16'h46F2;
 buffer[1798] = 16'h051E;
 buffer[1799] = 16'h0E04;
 buffer[1800] = 16'h2881;
 buffer[1801] = 16'h8029;
 buffer[1802] = 16'h46F2;
 buffer[1803] = 16'h0273;
 buffer[1804] = 16'h0E10;
 buffer[1805] = 16'h3C83;
 buffer[1806] = 16'h3E5C;
 buffer[1807] = 16'hFE86;
 buffer[1808] = 16'h6C00;
 buffer[1809] = 16'hFE84;
 buffer[1810] = 16'h6023;
 buffer[1811] = 16'h710F;
 buffer[1812] = 16'h0E1A;
 buffer[1813] = 16'h5C81;
 buffer[1814] = 16'hFEB6;
 buffer[1815] = 16'h03BC;
 buffer[1816] = 16'h0E2A;
 buffer[1817] = 16'h7704;
 buffer[1818] = 16'h726F;
 buffer[1819] = 16'h0064;
 buffer[1820] = 16'h46F2;
 buffer[1821] = 16'h4394;
 buffer[1822] = 16'h434B;
 buffer[1823] = 16'h05D3;
 buffer[1824] = 16'h0E32;
 buffer[1825] = 16'h7405;
 buffer[1826] = 16'h6B6F;
 buffer[1827] = 16'h6E65;
 buffer[1828] = 16'h435C;
 buffer[1829] = 16'h071C;
 buffer[1830] = 16'h0E42;
 buffer[1831] = 16'h6E05;
 buffer[1832] = 16'h6D61;
 buffer[1833] = 16'h3E65;
 buffer[1834] = 16'h438C;
 buffer[1835] = 16'h801F;
 buffer[1836] = 16'h6303;
 buffer[1837] = 16'h6203;
 buffer[1838] = 16'h039B;
 buffer[1839] = 16'h0E4E;
 buffer[1840] = 16'h7305;
 buffer[1841] = 16'h6D61;
 buffer[1842] = 16'h3F65;
 buffer[1843] = 16'h6A00;
 buffer[1844] = 16'h6147;
 buffer[1845] = 16'h0743;
 buffer[1846] = 16'h6181;
 buffer[1847] = 16'h6B81;
 buffer[1848] = 16'h6203;
 buffer[1849] = 16'h417E;
 buffer[1850] = 16'h6181;
 buffer[1851] = 16'h6B81;
 buffer[1852] = 16'h6203;
 buffer[1853] = 16'h417E;
 buffer[1854] = 16'h428F;
 buffer[1855] = 16'h4264;
 buffer[1856] = 16'h2743;
 buffer[1857] = 16'h6B8D;
 buffer[1858] = 16'h710F;
 buffer[1859] = 16'h6B81;
 buffer[1860] = 16'h2749;
 buffer[1861] = 16'h6B8D;
 buffer[1862] = 16'h6A00;
 buffer[1863] = 16'h6147;
 buffer[1864] = 16'h0736;
 buffer[1865] = 16'h6B8D;
 buffer[1866] = 16'h6103;
 buffer[1867] = 16'h8000;
 buffer[1868] = 16'h700C;
 buffer[1869] = 16'h0E60;
 buffer[1870] = 16'h6604;
 buffer[1871] = 16'h6E69;
 buffer[1872] = 16'h0064;
 buffer[1873] = 16'h6180;
 buffer[1874] = 16'h6081;
 buffer[1875] = 16'h417E;
 buffer[1876] = 16'hFE82;
 buffer[1877] = 16'h6023;
 buffer[1878] = 16'h6103;
 buffer[1879] = 16'h6081;
 buffer[1880] = 16'h6C00;
 buffer[1881] = 16'h6147;
 buffer[1882] = 16'h434B;
 buffer[1883] = 16'h6180;
 buffer[1884] = 16'h6C00;
 buffer[1885] = 16'h6081;
 buffer[1886] = 16'h276F;
 buffer[1887] = 16'h6081;
 buffer[1888] = 16'h6C00;
 buffer[1889] = 16'hFF1F;
 buffer[1890] = 16'h6303;
 buffer[1891] = 16'h6B81;
 buffer[1892] = 16'h6503;
 buffer[1893] = 16'h276A;
 buffer[1894] = 16'h434B;
 buffer[1895] = 16'h8000;
 buffer[1896] = 16'h6600;
 buffer[1897] = 16'h076E;
 buffer[1898] = 16'h434B;
 buffer[1899] = 16'hFE82;
 buffer[1900] = 16'h6C00;
 buffer[1901] = 16'h4733;
 buffer[1902] = 16'h0774;
 buffer[1903] = 16'h6B8D;
 buffer[1904] = 16'h6103;
 buffer[1905] = 16'h6180;
 buffer[1906] = 16'h4351;
 buffer[1907] = 16'h718C;
 buffer[1908] = 16'h2779;
 buffer[1909] = 16'h8002;
 buffer[1910] = 16'h4357;
 buffer[1911] = 16'h428F;
 buffer[1912] = 16'h075C;
 buffer[1913] = 16'h6B8D;
 buffer[1914] = 16'h6103;
 buffer[1915] = 16'h6003;
 buffer[1916] = 16'h4351;
 buffer[1917] = 16'h6081;
 buffer[1918] = 16'h472A;
 buffer[1919] = 16'h718C;
 buffer[1920] = 16'h0E9C;
 buffer[1921] = 16'h3C07;
 buffer[1922] = 16'h616E;
 buffer[1923] = 16'h656D;
 buffer[1924] = 16'h3E3F;
 buffer[1925] = 16'hFE90;
 buffer[1926] = 16'h6081;
 buffer[1927] = 16'h4383;
 buffer[1928] = 16'h6503;
 buffer[1929] = 16'h278B;
 buffer[1930] = 16'h4351;
 buffer[1931] = 16'h6147;
 buffer[1932] = 16'h6B8D;
 buffer[1933] = 16'h434B;
 buffer[1934] = 16'h6081;
 buffer[1935] = 16'h6147;
 buffer[1936] = 16'h6C00;
 buffer[1937] = 16'h4264;
 buffer[1938] = 16'h2798;
 buffer[1939] = 16'h4751;
 buffer[1940] = 16'h4264;
 buffer[1941] = 16'h278C;
 buffer[1942] = 16'h6B8D;
 buffer[1943] = 16'h710F;
 buffer[1944] = 16'h6B8D;
 buffer[1945] = 16'h6103;
 buffer[1946] = 16'h8000;
 buffer[1947] = 16'h700C;
 buffer[1948] = 16'h0F02;
 buffer[1949] = 16'h6E05;
 buffer[1950] = 16'h6D61;
 buffer[1951] = 16'h3F65;
 buffer[1952] = 16'hFEB8;
 buffer[1953] = 16'h03BC;
 buffer[1954] = 16'h0F3A;
 buffer[1955] = 16'h5E02;
 buffer[1956] = 16'h0068;
 buffer[1957] = 16'h6147;
 buffer[1958] = 16'h6181;
 buffer[1959] = 16'h6B81;
 buffer[1960] = 16'h6803;
 buffer[1961] = 16'h6081;
 buffer[1962] = 16'h27B0;
 buffer[1963] = 16'h8008;
 buffer[1964] = 16'h6081;
 buffer[1965] = 16'h44CC;
 buffer[1966] = 16'h4506;
 buffer[1967] = 16'h44CC;
 buffer[1968] = 16'h6B8D;
 buffer[1969] = 16'h720F;
 buffer[1970] = 16'h0F46;
 buffer[1971] = 16'h7403;
 buffer[1972] = 16'h7061;
 buffer[1973] = 16'h6081;
 buffer[1974] = 16'h44CC;
 buffer[1975] = 16'h6181;
 buffer[1976] = 16'h418D;
 buffer[1977] = 16'h731C;
 buffer[1978] = 16'h0F66;
 buffer[1979] = 16'h6B04;
 buffer[1980] = 16'h6174;
 buffer[1981] = 16'h0070;
 buffer[1982] = 16'h6081;
 buffer[1983] = 16'h800D;
 buffer[1984] = 16'h6503;
 buffer[1985] = 16'h27C8;
 buffer[1986] = 16'h8008;
 buffer[1987] = 16'h6503;
 buffer[1988] = 16'h27C7;
 buffer[1989] = 16'h435C;
 buffer[1990] = 16'h07B5;
 buffer[1991] = 16'h07A5;
 buffer[1992] = 16'h6103;
 buffer[1993] = 16'h6003;
 buffer[1994] = 16'h708D;
 buffer[1995] = 16'h0F76;
 buffer[1996] = 16'h6106;
 buffer[1997] = 16'h6363;
 buffer[1998] = 16'h7065;
 buffer[1999] = 16'h0074;
 buffer[2000] = 16'h6181;
 buffer[2001] = 16'h6203;
 buffer[2002] = 16'h6181;
 buffer[2003] = 16'h4279;
 buffer[2004] = 16'h6503;
 buffer[2005] = 16'h27E1;
 buffer[2006] = 16'h44D1;
 buffer[2007] = 16'h6081;
 buffer[2008] = 16'h435C;
 buffer[2009] = 16'h428F;
 buffer[2010] = 16'h807F;
 buffer[2011] = 16'h6F03;
 buffer[2012] = 16'h27DF;
 buffer[2013] = 16'h47B5;
 buffer[2014] = 16'h07E0;
 buffer[2015] = 16'h47BE;
 buffer[2016] = 16'h07D3;
 buffer[2017] = 16'h6103;
 buffer[2018] = 16'h6181;
 buffer[2019] = 16'h028F;
 buffer[2020] = 16'h0F98;
 buffer[2021] = 16'h7105;
 buffer[2022] = 16'h6575;
 buffer[2023] = 16'h7972;
 buffer[2024] = 16'hFE88;
 buffer[2025] = 16'h6C00;
 buffer[2026] = 16'h8050;
 buffer[2027] = 16'h47D0;
 buffer[2028] = 16'hFE86;
 buffer[2029] = 16'h6023;
 buffer[2030] = 16'h6103;
 buffer[2031] = 16'h6103;
 buffer[2032] = 16'h8000;
 buffer[2033] = 16'hFE84;
 buffer[2034] = 16'h6023;
 buffer[2035] = 16'h710F;
 buffer[2036] = 16'h0FCA;
 buffer[2037] = 16'h6106;
 buffer[2038] = 16'h6F62;
 buffer[2039] = 16'h7472;
 buffer[2040] = 16'h0032;
 buffer[2041] = 16'h4535;
 buffer[2042] = 16'h710F;
 buffer[2043] = 16'h0FEA;
 buffer[2044] = 16'h6106;
 buffer[2045] = 16'h6F62;
 buffer[2046] = 16'h7472;
 buffer[2047] = 16'h0031;
 buffer[2048] = 16'h4506;
 buffer[2049] = 16'h4547;
 buffer[2050] = 16'h803F;
 buffer[2051] = 16'h44CC;
 buffer[2052] = 16'h452E;
 buffer[2053] = 16'hFE8C;
 buffer[2054] = 16'h43BC;
 buffer[2055] = 16'h07F9;
 buffer[2056] = 16'h0FF8;
 buffer[2057] = 16'h3C49;
 buffer[2058] = 16'h613F;
 buffer[2059] = 16'h6F62;
 buffer[2060] = 16'h7472;
 buffer[2061] = 16'h3E22;
 buffer[2062] = 16'h2811;
 buffer[2063] = 16'h4535;
 buffer[2064] = 16'h0800;
 buffer[2065] = 16'h07F9;
 buffer[2066] = 16'h1012;
 buffer[2067] = 16'h6606;
 buffer[2068] = 16'h726F;
 buffer[2069] = 16'h6567;
 buffer[2070] = 16'h0074;
 buffer[2071] = 16'h4724;
 buffer[2072] = 16'h47A0;
 buffer[2073] = 16'h4264;
 buffer[2074] = 16'h2829;
 buffer[2075] = 16'h4351;
 buffer[2076] = 16'h6081;
 buffer[2077] = 16'hFEAC;
 buffer[2078] = 16'h6023;
 buffer[2079] = 16'h6103;
 buffer[2080] = 16'h6C00;
 buffer[2081] = 16'h6081;
 buffer[2082] = 16'hFE90;
 buffer[2083] = 16'h6023;
 buffer[2084] = 16'h6103;
 buffer[2085] = 16'hFEAE;
 buffer[2086] = 16'h6023;
 buffer[2087] = 16'h6103;
 buffer[2088] = 16'h710F;
 buffer[2089] = 16'h0800;
 buffer[2090] = 16'h1026;
 buffer[2091] = 16'h240A;
 buffer[2092] = 16'h6E69;
 buffer[2093] = 16'h6574;
 buffer[2094] = 16'h7072;
 buffer[2095] = 16'h6572;
 buffer[2096] = 16'h0074;
 buffer[2097] = 16'h47A0;
 buffer[2098] = 16'h4264;
 buffer[2099] = 16'h2841;
 buffer[2100] = 16'h6C00;
 buffer[2101] = 16'h8040;
 buffer[2102] = 16'h6303;
 buffer[2103] = 16'h480E;
 buffer[2104] = 16'h630C;
 buffer[2105] = 16'h6D6F;
 buffer[2106] = 16'h6970;
 buffer[2107] = 16'h656C;
 buffer[2108] = 16'h6F2D;
 buffer[2109] = 16'h6C6E;
 buffer[2110] = 16'h0079;
 buffer[2111] = 16'h0172;
 buffer[2112] = 16'h0845;
 buffer[2113] = 16'h445F;
 buffer[2114] = 16'h2844;
 buffer[2115] = 16'h700C;
 buffer[2116] = 16'h0800;
 buffer[2117] = 16'h1056;
 buffer[2118] = 16'h5B81;
 buffer[2119] = 16'h9062;
 buffer[2120] = 16'hFE8A;
 buffer[2121] = 16'h6023;
 buffer[2122] = 16'h710F;
 buffer[2123] = 16'h108C;
 buffer[2124] = 16'h2E03;
 buffer[2125] = 16'h6B6F;
 buffer[2126] = 16'h9062;
 buffer[2127] = 16'hFE8A;
 buffer[2128] = 16'h6C00;
 buffer[2129] = 16'h6703;
 buffer[2130] = 16'h2856;
 buffer[2131] = 16'h454C;
 buffer[2132] = 16'h2003;
 buffer[2133] = 16'h6B6F;
 buffer[2134] = 16'h052E;
 buffer[2135] = 16'h1098;
 buffer[2136] = 16'h6504;
 buffer[2137] = 16'h6176;
 buffer[2138] = 16'h006C;
 buffer[2139] = 16'h4724;
 buffer[2140] = 16'h6081;
 buffer[2141] = 16'h417E;
 buffer[2142] = 16'h2862;
 buffer[2143] = 16'hFE8A;
 buffer[2144] = 16'h43BC;
 buffer[2145] = 16'h085B;
 buffer[2146] = 16'h6103;
 buffer[2147] = 16'h084E;
 buffer[2148] = 16'h10B0;
 buffer[2149] = 16'h2445;
 buffer[2150] = 16'h7665;
 buffer[2151] = 16'h6C61;
 buffer[2152] = 16'hFE84;
 buffer[2153] = 16'h6C00;
 buffer[2154] = 16'h6147;
 buffer[2155] = 16'hFE86;
 buffer[2156] = 16'h6C00;
 buffer[2157] = 16'h6147;
 buffer[2158] = 16'hFE88;
 buffer[2159] = 16'h6C00;
 buffer[2160] = 16'h6147;
 buffer[2161] = 16'hFE84;
 buffer[2162] = 16'h8000;
 buffer[2163] = 16'h6180;
 buffer[2164] = 16'h6023;
 buffer[2165] = 16'h6103;
 buffer[2166] = 16'hFE86;
 buffer[2167] = 16'h6023;
 buffer[2168] = 16'h6103;
 buffer[2169] = 16'hFE88;
 buffer[2170] = 16'h6023;
 buffer[2171] = 16'h6103;
 buffer[2172] = 16'h485B;
 buffer[2173] = 16'h6B8D;
 buffer[2174] = 16'hFE88;
 buffer[2175] = 16'h6023;
 buffer[2176] = 16'h6103;
 buffer[2177] = 16'h6B8D;
 buffer[2178] = 16'hFE86;
 buffer[2179] = 16'h6023;
 buffer[2180] = 16'h6103;
 buffer[2181] = 16'h6B8D;
 buffer[2182] = 16'hFE84;
 buffer[2183] = 16'h6023;
 buffer[2184] = 16'h710F;
 buffer[2185] = 16'h10CA;
 buffer[2186] = 16'h7006;
 buffer[2187] = 16'h6572;
 buffer[2188] = 16'h6573;
 buffer[2189] = 16'h0074;
 buffer[2190] = 16'hFF00;
 buffer[2191] = 16'hFE86;
 buffer[2192] = 16'h434B;
 buffer[2193] = 16'h6023;
 buffer[2194] = 16'h710F;
 buffer[2195] = 16'h1114;
 buffer[2196] = 16'h7104;
 buffer[2197] = 16'h6975;
 buffer[2198] = 16'h0074;
 buffer[2199] = 16'h4847;
 buffer[2200] = 16'h47E8;
 buffer[2201] = 16'h485B;
 buffer[2202] = 16'h0898;
 buffer[2203] = 16'h700C;
 buffer[2204] = 16'h1128;
 buffer[2205] = 16'h6105;
 buffer[2206] = 16'h6F62;
 buffer[2207] = 16'h7472;
 buffer[2208] = 16'h6103;
 buffer[2209] = 16'h488E;
 buffer[2210] = 16'h484E;
 buffer[2211] = 16'h0897;
 buffer[2212] = 16'h113A;
 buffer[2213] = 16'h2701;
 buffer[2214] = 16'h4724;
 buffer[2215] = 16'h47A0;
 buffer[2216] = 16'h28AA;
 buffer[2217] = 16'h700C;
 buffer[2218] = 16'h0800;
 buffer[2219] = 16'h114A;
 buffer[2220] = 16'h6105;
 buffer[2221] = 16'h6C6C;
 buffer[2222] = 16'h746F;
 buffer[2223] = 16'h439B;
 buffer[2224] = 16'hFEAC;
 buffer[2225] = 16'h0370;
 buffer[2226] = 16'h1158;
 buffer[2227] = 16'h2C01;
 buffer[2228] = 16'h4394;
 buffer[2229] = 16'h6081;
 buffer[2230] = 16'h434B;
 buffer[2231] = 16'hFEAC;
 buffer[2232] = 16'h6023;
 buffer[2233] = 16'h6103;
 buffer[2234] = 16'h6023;
 buffer[2235] = 16'h710F;
 buffer[2236] = 16'h1166;
 buffer[2237] = 16'h6345;
 buffer[2238] = 16'h6C61;
 buffer[2239] = 16'h2C6C;
 buffer[2240] = 16'h8001;
 buffer[2241] = 16'h6903;
 buffer[2242] = 16'hC000;
 buffer[2243] = 16'h6403;
 buffer[2244] = 16'h08B4;
 buffer[2245] = 16'h117A;
 buffer[2246] = 16'h3F47;
 buffer[2247] = 16'h7262;
 buffer[2248] = 16'h6E61;
 buffer[2249] = 16'h6863;
 buffer[2250] = 16'h8001;
 buffer[2251] = 16'h6903;
 buffer[2252] = 16'hA000;
 buffer[2253] = 16'h6403;
 buffer[2254] = 16'h08B4;
 buffer[2255] = 16'h118C;
 buffer[2256] = 16'h6246;
 buffer[2257] = 16'h6172;
 buffer[2258] = 16'h636E;
 buffer[2259] = 16'h0068;
 buffer[2260] = 16'h8001;
 buffer[2261] = 16'h6903;
 buffer[2262] = 16'h8000;
 buffer[2263] = 16'h6403;
 buffer[2264] = 16'h08B4;
 buffer[2265] = 16'h11A0;
 buffer[2266] = 16'h5B89;
 buffer[2267] = 16'h6F63;
 buffer[2268] = 16'h706D;
 buffer[2269] = 16'h6C69;
 buffer[2270] = 16'h5D65;
 buffer[2271] = 16'h48A6;
 buffer[2272] = 16'h08C0;
 buffer[2273] = 16'h11B4;
 buffer[2274] = 16'h6347;
 buffer[2275] = 16'h6D6F;
 buffer[2276] = 16'h6970;
 buffer[2277] = 16'h656C;
 buffer[2278] = 16'h6B8D;
 buffer[2279] = 16'h6081;
 buffer[2280] = 16'h6C00;
 buffer[2281] = 16'h48B4;
 buffer[2282] = 16'h434B;
 buffer[2283] = 16'h6147;
 buffer[2284] = 16'h700C;
 buffer[2285] = 16'h11C4;
 buffer[2286] = 16'h7287;
 buffer[2287] = 16'h6365;
 buffer[2288] = 16'h7275;
 buffer[2289] = 16'h6573;
 buffer[2290] = 16'hFEAE;
 buffer[2291] = 16'h6C00;
 buffer[2292] = 16'h472A;
 buffer[2293] = 16'h08C0;
 buffer[2294] = 16'h11DC;
 buffer[2295] = 16'h7004;
 buffer[2296] = 16'h6369;
 buffer[2297] = 16'h006B;
 buffer[2298] = 16'h6081;
 buffer[2299] = 16'h6410;
 buffer[2300] = 16'h6410;
 buffer[2301] = 16'h80C0;
 buffer[2302] = 16'h6203;
 buffer[2303] = 16'h6147;
 buffer[2304] = 16'h700C;
 buffer[2305] = 16'h11EE;
 buffer[2306] = 16'h6C87;
 buffer[2307] = 16'h7469;
 buffer[2308] = 16'h7265;
 buffer[2309] = 16'h6C61;
 buffer[2310] = 16'h6081;
 buffer[2311] = 16'hFFFF;
 buffer[2312] = 16'h6600;
 buffer[2313] = 16'h6303;
 buffer[2314] = 16'h2912;
 buffer[2315] = 16'h8000;
 buffer[2316] = 16'h6600;
 buffer[2317] = 16'h6503;
 buffer[2318] = 16'h4906;
 buffer[2319] = 16'h48E6;
 buffer[2320] = 16'h6600;
 buffer[2321] = 16'h0916;
 buffer[2322] = 16'hFFFF;
 buffer[2323] = 16'h6600;
 buffer[2324] = 16'h6403;
 buffer[2325] = 16'h08B4;
 buffer[2326] = 16'h700C;
 buffer[2327] = 16'h1204;
 buffer[2328] = 16'h5B83;
 buffer[2329] = 16'h5D27;
 buffer[2330] = 16'h48A6;
 buffer[2331] = 16'h0906;
 buffer[2332] = 16'h1230;
 buffer[2333] = 16'h2403;
 buffer[2334] = 16'h222C;
 buffer[2335] = 16'h8022;
 buffer[2336] = 16'h46F2;
 buffer[2337] = 16'h4394;
 buffer[2338] = 16'h45D3;
 buffer[2339] = 16'h438C;
 buffer[2340] = 16'h6203;
 buffer[2341] = 16'h439B;
 buffer[2342] = 16'hFEAC;
 buffer[2343] = 16'h6023;
 buffer[2344] = 16'h710F;
 buffer[2345] = 16'h123A;
 buffer[2346] = 16'h66C3;
 buffer[2347] = 16'h726F;
 buffer[2348] = 16'h48E6;
 buffer[2349] = 16'h4112;
 buffer[2350] = 16'h0394;
 buffer[2351] = 16'h1254;
 buffer[2352] = 16'h62C5;
 buffer[2353] = 16'h6765;
 buffer[2354] = 16'h6E69;
 buffer[2355] = 16'h0394;
 buffer[2356] = 16'h1260;
 buffer[2357] = 16'h2846;
 buffer[2358] = 16'h656E;
 buffer[2359] = 16'h7478;
 buffer[2360] = 16'h0029;
 buffer[2361] = 16'h6B8D;
 buffer[2362] = 16'h6B8D;
 buffer[2363] = 16'h4264;
 buffer[2364] = 16'h2942;
 buffer[2365] = 16'h6A00;
 buffer[2366] = 16'h6147;
 buffer[2367] = 16'h6C00;
 buffer[2368] = 16'h6147;
 buffer[2369] = 16'h700C;
 buffer[2370] = 16'h434B;
 buffer[2371] = 16'h6147;
 buffer[2372] = 16'h700C;
 buffer[2373] = 16'h126A;
 buffer[2374] = 16'h6EC4;
 buffer[2375] = 16'h7865;
 buffer[2376] = 16'h0074;
 buffer[2377] = 16'h48E6;
 buffer[2378] = 16'h4939;
 buffer[2379] = 16'h08B4;
 buffer[2380] = 16'h128C;
 buffer[2381] = 16'h2844;
 buffer[2382] = 16'h6F64;
 buffer[2383] = 16'h0029;
 buffer[2384] = 16'h6B8D;
 buffer[2385] = 16'h6081;
 buffer[2386] = 16'h6147;
 buffer[2387] = 16'h6180;
 buffer[2388] = 16'h426B;
 buffer[2389] = 16'h6147;
 buffer[2390] = 16'h6147;
 buffer[2391] = 16'h434B;
 buffer[2392] = 16'h6147;
 buffer[2393] = 16'h700C;
 buffer[2394] = 16'h129A;
 buffer[2395] = 16'h64C2;
 buffer[2396] = 16'h006F;
 buffer[2397] = 16'h48E6;
 buffer[2398] = 16'h4950;
 buffer[2399] = 16'h8000;
 buffer[2400] = 16'h48B4;
 buffer[2401] = 16'h0394;
 buffer[2402] = 16'h12B6;
 buffer[2403] = 16'h2847;
 buffer[2404] = 16'h656C;
 buffer[2405] = 16'h7661;
 buffer[2406] = 16'h2965;
 buffer[2407] = 16'h6B8D;
 buffer[2408] = 16'h6103;
 buffer[2409] = 16'h6B8D;
 buffer[2410] = 16'h6103;
 buffer[2411] = 16'h6B8D;
 buffer[2412] = 16'h710F;
 buffer[2413] = 16'h12C6;
 buffer[2414] = 16'h6CC5;
 buffer[2415] = 16'h6165;
 buffer[2416] = 16'h6576;
 buffer[2417] = 16'h48E6;
 buffer[2418] = 16'h4967;
 buffer[2419] = 16'h700C;
 buffer[2420] = 16'h12DC;
 buffer[2421] = 16'h2846;
 buffer[2422] = 16'h6F6C;
 buffer[2423] = 16'h706F;
 buffer[2424] = 16'h0029;
 buffer[2425] = 16'h6B8D;
 buffer[2426] = 16'h6B8D;
 buffer[2427] = 16'h6310;
 buffer[2428] = 16'h6B8D;
 buffer[2429] = 16'h4279;
 buffer[2430] = 16'h6213;
 buffer[2431] = 16'h2985;
 buffer[2432] = 16'h6147;
 buffer[2433] = 16'h6147;
 buffer[2434] = 16'h6C00;
 buffer[2435] = 16'h6147;
 buffer[2436] = 16'h700C;
 buffer[2437] = 16'h6147;
 buffer[2438] = 16'h6A00;
 buffer[2439] = 16'h6147;
 buffer[2440] = 16'h434B;
 buffer[2441] = 16'h6147;
 buffer[2442] = 16'h700C;
 buffer[2443] = 16'h12EA;
 buffer[2444] = 16'h2848;
 buffer[2445] = 16'h6E75;
 buffer[2446] = 16'h6F6C;
 buffer[2447] = 16'h706F;
 buffer[2448] = 16'h0029;
 buffer[2449] = 16'h6B8D;
 buffer[2450] = 16'h6B8D;
 buffer[2451] = 16'h6103;
 buffer[2452] = 16'h6B8D;
 buffer[2453] = 16'h6103;
 buffer[2454] = 16'h6B8D;
 buffer[2455] = 16'h6103;
 buffer[2456] = 16'h6147;
 buffer[2457] = 16'h700C;
 buffer[2458] = 16'h1318;
 buffer[2459] = 16'h75C6;
 buffer[2460] = 16'h6C6E;
 buffer[2461] = 16'h6F6F;
 buffer[2462] = 16'h0070;
 buffer[2463] = 16'h48E6;
 buffer[2464] = 16'h4991;
 buffer[2465] = 16'h700C;
 buffer[2466] = 16'h1336;
 buffer[2467] = 16'h2845;
 buffer[2468] = 16'h643F;
 buffer[2469] = 16'h296F;
 buffer[2470] = 16'h4279;
 buffer[2471] = 16'h6213;
 buffer[2472] = 16'h29B3;
 buffer[2473] = 16'h6B8D;
 buffer[2474] = 16'h6081;
 buffer[2475] = 16'h6147;
 buffer[2476] = 16'h6180;
 buffer[2477] = 16'h426B;
 buffer[2478] = 16'h6147;
 buffer[2479] = 16'h6147;
 buffer[2480] = 16'h434B;
 buffer[2481] = 16'h6147;
 buffer[2482] = 16'h700C;
 buffer[2483] = 16'h0273;
 buffer[2484] = 16'h700C;
 buffer[2485] = 16'h1346;
 buffer[2486] = 16'h3FC3;
 buffer[2487] = 16'h6F64;
 buffer[2488] = 16'h48E6;
 buffer[2489] = 16'h49A6;
 buffer[2490] = 16'h8000;
 buffer[2491] = 16'h48B4;
 buffer[2492] = 16'h0394;
 buffer[2493] = 16'h136C;
 buffer[2494] = 16'h6CC4;
 buffer[2495] = 16'h6F6F;
 buffer[2496] = 16'h0070;
 buffer[2497] = 16'h48E6;
 buffer[2498] = 16'h4979;
 buffer[2499] = 16'h6081;
 buffer[2500] = 16'h48B4;
 buffer[2501] = 16'h48E6;
 buffer[2502] = 16'h4991;
 buffer[2503] = 16'h4351;
 buffer[2504] = 16'h4394;
 buffer[2505] = 16'h8001;
 buffer[2506] = 16'h6903;
 buffer[2507] = 16'h6180;
 buffer[2508] = 16'h6023;
 buffer[2509] = 16'h710F;
 buffer[2510] = 16'h137C;
 buffer[2511] = 16'h2847;
 buffer[2512] = 16'h6C2B;
 buffer[2513] = 16'h6F6F;
 buffer[2514] = 16'h2970;
 buffer[2515] = 16'h6B8D;
 buffer[2516] = 16'h6180;
 buffer[2517] = 16'h6B8D;
 buffer[2518] = 16'h6B8D;
 buffer[2519] = 16'h4279;
 buffer[2520] = 16'h428F;
 buffer[2521] = 16'h6147;
 buffer[2522] = 16'h8002;
 buffer[2523] = 16'h48FA;
 buffer[2524] = 16'h6B81;
 buffer[2525] = 16'h6203;
 buffer[2526] = 16'h6B81;
 buffer[2527] = 16'h6503;
 buffer[2528] = 16'h6810;
 buffer[2529] = 16'h6010;
 buffer[2530] = 16'h8003;
 buffer[2531] = 16'h48FA;
 buffer[2532] = 16'h6B8D;
 buffer[2533] = 16'h6503;
 buffer[2534] = 16'h6810;
 buffer[2535] = 16'h6010;
 buffer[2536] = 16'h6403;
 buffer[2537] = 16'h29F0;
 buffer[2538] = 16'h6147;
 buffer[2539] = 16'h6203;
 buffer[2540] = 16'h6147;
 buffer[2541] = 16'h6C00;
 buffer[2542] = 16'h6147;
 buffer[2543] = 16'h700C;
 buffer[2544] = 16'h6147;
 buffer[2545] = 16'h6147;
 buffer[2546] = 16'h6103;
 buffer[2547] = 16'h434B;
 buffer[2548] = 16'h6147;
 buffer[2549] = 16'h700C;
 buffer[2550] = 16'h139E;
 buffer[2551] = 16'h2BC5;
 buffer[2552] = 16'h6F6C;
 buffer[2553] = 16'h706F;
 buffer[2554] = 16'h48E6;
 buffer[2555] = 16'h49D3;
 buffer[2556] = 16'h6081;
 buffer[2557] = 16'h48B4;
 buffer[2558] = 16'h48E6;
 buffer[2559] = 16'h4991;
 buffer[2560] = 16'h4351;
 buffer[2561] = 16'h4394;
 buffer[2562] = 16'h8001;
 buffer[2563] = 16'h6903;
 buffer[2564] = 16'h6180;
 buffer[2565] = 16'h6023;
 buffer[2566] = 16'h710F;
 buffer[2567] = 16'h13EE;
 buffer[2568] = 16'h2843;
 buffer[2569] = 16'h2969;
 buffer[2570] = 16'h6B8D;
 buffer[2571] = 16'h6B8D;
 buffer[2572] = 16'h414F;
 buffer[2573] = 16'h6147;
 buffer[2574] = 16'h6147;
 buffer[2575] = 16'h700C;
 buffer[2576] = 16'h1410;
 buffer[2577] = 16'h69C1;
 buffer[2578] = 16'h48E6;
 buffer[2579] = 16'h4A0A;
 buffer[2580] = 16'h700C;
 buffer[2581] = 16'h1422;
 buffer[2582] = 16'h75C5;
 buffer[2583] = 16'h746E;
 buffer[2584] = 16'h6C69;
 buffer[2585] = 16'h08CA;
 buffer[2586] = 16'h142C;
 buffer[2587] = 16'h61C5;
 buffer[2588] = 16'h6167;
 buffer[2589] = 16'h6E69;
 buffer[2590] = 16'h08D4;
 buffer[2591] = 16'h1436;
 buffer[2592] = 16'h69C2;
 buffer[2593] = 16'h0066;
 buffer[2594] = 16'h4394;
 buffer[2595] = 16'h8000;
 buffer[2596] = 16'h08CA;
 buffer[2597] = 16'h1440;
 buffer[2598] = 16'h74C4;
 buffer[2599] = 16'h6568;
 buffer[2600] = 16'h006E;
 buffer[2601] = 16'h4394;
 buffer[2602] = 16'h8001;
 buffer[2603] = 16'h6903;
 buffer[2604] = 16'h6181;
 buffer[2605] = 16'h6C00;
 buffer[2606] = 16'h6403;
 buffer[2607] = 16'h6180;
 buffer[2608] = 16'h6023;
 buffer[2609] = 16'h710F;
 buffer[2610] = 16'h144C;
 buffer[2611] = 16'h72C6;
 buffer[2612] = 16'h7065;
 buffer[2613] = 16'h6165;
 buffer[2614] = 16'h0074;
 buffer[2615] = 16'h48D4;
 buffer[2616] = 16'h0A29;
 buffer[2617] = 16'h1466;
 buffer[2618] = 16'h73C4;
 buffer[2619] = 16'h696B;
 buffer[2620] = 16'h0070;
 buffer[2621] = 16'h4394;
 buffer[2622] = 16'h8000;
 buffer[2623] = 16'h08D4;
 buffer[2624] = 16'h1474;
 buffer[2625] = 16'h61C3;
 buffer[2626] = 16'h7466;
 buffer[2627] = 16'h6103;
 buffer[2628] = 16'h4A3D;
 buffer[2629] = 16'h4933;
 buffer[2630] = 16'h718C;
 buffer[2631] = 16'h1482;
 buffer[2632] = 16'h65C4;
 buffer[2633] = 16'h736C;
 buffer[2634] = 16'h0065;
 buffer[2635] = 16'h4A3D;
 buffer[2636] = 16'h6180;
 buffer[2637] = 16'h0A29;
 buffer[2638] = 16'h1490;
 buffer[2639] = 16'h77C5;
 buffer[2640] = 16'h6968;
 buffer[2641] = 16'h656C;
 buffer[2642] = 16'h4A22;
 buffer[2643] = 16'h718C;
 buffer[2644] = 16'h149E;
 buffer[2645] = 16'h2846;
 buffer[2646] = 16'h6163;
 buffer[2647] = 16'h6573;
 buffer[2648] = 16'h0029;
 buffer[2649] = 16'h6B8D;
 buffer[2650] = 16'h6180;
 buffer[2651] = 16'h6147;
 buffer[2652] = 16'h6147;
 buffer[2653] = 16'h700C;
 buffer[2654] = 16'h14AA;
 buffer[2655] = 16'h63C4;
 buffer[2656] = 16'h7361;
 buffer[2657] = 16'h0065;
 buffer[2658] = 16'h48E6;
 buffer[2659] = 16'h4A59;
 buffer[2660] = 16'h8030;
 buffer[2661] = 16'h700C;
 buffer[2662] = 16'h14BE;
 buffer[2663] = 16'h2844;
 buffer[2664] = 16'h666F;
 buffer[2665] = 16'h0029;
 buffer[2666] = 16'h6B8D;
 buffer[2667] = 16'h6B81;
 buffer[2668] = 16'h6180;
 buffer[2669] = 16'h6147;
 buffer[2670] = 16'h770F;
 buffer[2671] = 16'h14CE;
 buffer[2672] = 16'h6FC2;
 buffer[2673] = 16'h0066;
 buffer[2674] = 16'h48E6;
 buffer[2675] = 16'h4A6A;
 buffer[2676] = 16'h0A22;
 buffer[2677] = 16'h14E0;
 buffer[2678] = 16'h65C5;
 buffer[2679] = 16'h646E;
 buffer[2680] = 16'h666F;
 buffer[2681] = 16'h4A4B;
 buffer[2682] = 16'h8031;
 buffer[2683] = 16'h700C;
 buffer[2684] = 16'h14EC;
 buffer[2685] = 16'h2809;
 buffer[2686] = 16'h6E65;
 buffer[2687] = 16'h6364;
 buffer[2688] = 16'h7361;
 buffer[2689] = 16'h2965;
 buffer[2690] = 16'h6B8D;
 buffer[2691] = 16'h6B8D;
 buffer[2692] = 16'h6103;
 buffer[2693] = 16'h6147;
 buffer[2694] = 16'h700C;
 buffer[2695] = 16'h14FA;
 buffer[2696] = 16'h65C7;
 buffer[2697] = 16'h646E;
 buffer[2698] = 16'h6163;
 buffer[2699] = 16'h6573;
 buffer[2700] = 16'h6081;
 buffer[2701] = 16'h8031;
 buffer[2702] = 16'h6703;
 buffer[2703] = 16'h2A93;
 buffer[2704] = 16'h6103;
 buffer[2705] = 16'h4A29;
 buffer[2706] = 16'h0A8C;
 buffer[2707] = 16'h8030;
 buffer[2708] = 16'h6213;
 buffer[2709] = 16'h480E;
 buffer[2710] = 16'h6213;
 buffer[2711] = 16'h6461;
 buffer[2712] = 16'h6320;
 buffer[2713] = 16'h7361;
 buffer[2714] = 16'h2065;
 buffer[2715] = 16'h6F63;
 buffer[2716] = 16'h736E;
 buffer[2717] = 16'h7274;
 buffer[2718] = 16'h6375;
 buffer[2719] = 16'h2E74;
 buffer[2720] = 16'h48E6;
 buffer[2721] = 16'h4A82;
 buffer[2722] = 16'h700C;
 buffer[2723] = 16'h1510;
 buffer[2724] = 16'h24C2;
 buffer[2725] = 16'h0022;
 buffer[2726] = 16'h48E6;
 buffer[2727] = 16'h4542;
 buffer[2728] = 16'h091F;
 buffer[2729] = 16'h1548;
 buffer[2730] = 16'h2EC2;
 buffer[2731] = 16'h0022;
 buffer[2732] = 16'h48E6;
 buffer[2733] = 16'h454C;
 buffer[2734] = 16'h091F;
 buffer[2735] = 16'h1554;
 buffer[2736] = 16'h3E05;
 buffer[2737] = 16'h6F62;
 buffer[2738] = 16'h7964;
 buffer[2739] = 16'h034B;
 buffer[2740] = 16'h1560;
 buffer[2741] = 16'h2844;
 buffer[2742] = 16'h6F74;
 buffer[2743] = 16'h0029;
 buffer[2744] = 16'h6B8D;
 buffer[2745] = 16'h6081;
 buffer[2746] = 16'h434B;
 buffer[2747] = 16'h6147;
 buffer[2748] = 16'h6C00;
 buffer[2749] = 16'h6023;
 buffer[2750] = 16'h710F;
 buffer[2751] = 16'h156A;
 buffer[2752] = 16'h74C2;
 buffer[2753] = 16'h006F;
 buffer[2754] = 16'h48E6;
 buffer[2755] = 16'h4AB8;
 buffer[2756] = 16'h48A6;
 buffer[2757] = 16'h4AB3;
 buffer[2758] = 16'h08B4;
 buffer[2759] = 16'h1580;
 buffer[2760] = 16'h2845;
 buffer[2761] = 16'h742B;
 buffer[2762] = 16'h296F;
 buffer[2763] = 16'h6B8D;
 buffer[2764] = 16'h6081;
 buffer[2765] = 16'h434B;
 buffer[2766] = 16'h6147;
 buffer[2767] = 16'h6C00;
 buffer[2768] = 16'h0370;
 buffer[2769] = 16'h1590;
 buffer[2770] = 16'h2BC3;
 buffer[2771] = 16'h6F74;
 buffer[2772] = 16'h48E6;
 buffer[2773] = 16'h4ACB;
 buffer[2774] = 16'h48A6;
 buffer[2775] = 16'h4AB3;
 buffer[2776] = 16'h08B4;
 buffer[2777] = 16'h15A4;
 buffer[2778] = 16'h670B;
 buffer[2779] = 16'h7465;
 buffer[2780] = 16'h632D;
 buffer[2781] = 16'h7275;
 buffer[2782] = 16'h6572;
 buffer[2783] = 16'h746E;
 buffer[2784] = 16'hFEA8;
 buffer[2785] = 16'h7C0C;
 buffer[2786] = 16'h15B4;
 buffer[2787] = 16'h730B;
 buffer[2788] = 16'h7465;
 buffer[2789] = 16'h632D;
 buffer[2790] = 16'h7275;
 buffer[2791] = 16'h6572;
 buffer[2792] = 16'h746E;
 buffer[2793] = 16'hFEA8;
 buffer[2794] = 16'h6023;
 buffer[2795] = 16'h710F;
 buffer[2796] = 16'h15C6;
 buffer[2797] = 16'h640B;
 buffer[2798] = 16'h6665;
 buffer[2799] = 16'h6E69;
 buffer[2800] = 16'h7469;
 buffer[2801] = 16'h6F69;
 buffer[2802] = 16'h736E;
 buffer[2803] = 16'hFE90;
 buffer[2804] = 16'h6C00;
 buffer[2805] = 16'h0AE9;
 buffer[2806] = 16'h15DA;
 buffer[2807] = 16'h3F07;
 buffer[2808] = 16'h6E75;
 buffer[2809] = 16'h7169;
 buffer[2810] = 16'h6575;
 buffer[2811] = 16'h6081;
 buffer[2812] = 16'h4AE0;
 buffer[2813] = 16'h4751;
 buffer[2814] = 16'h2B06;
 buffer[2815] = 16'h454C;
 buffer[2816] = 16'h2007;
 buffer[2817] = 16'h6572;
 buffer[2818] = 16'h6564;
 buffer[2819] = 16'h2066;
 buffer[2820] = 16'h6181;
 buffer[2821] = 16'h4547;
 buffer[2822] = 16'h710F;
 buffer[2823] = 16'h15EE;
 buffer[2824] = 16'h3C05;
 buffer[2825] = 16'h2C24;
 buffer[2826] = 16'h3E6E;
 buffer[2827] = 16'h6081;
 buffer[2828] = 16'h417E;
 buffer[2829] = 16'h2B20;
 buffer[2830] = 16'h4AFB;
 buffer[2831] = 16'h6081;
 buffer[2832] = 16'h438C;
 buffer[2833] = 16'h6203;
 buffer[2834] = 16'h439B;
 buffer[2835] = 16'hFEAC;
 buffer[2836] = 16'h6023;
 buffer[2837] = 16'h6103;
 buffer[2838] = 16'h6081;
 buffer[2839] = 16'hFEAE;
 buffer[2840] = 16'h6023;
 buffer[2841] = 16'h6103;
 buffer[2842] = 16'h4351;
 buffer[2843] = 16'h4AE0;
 buffer[2844] = 16'h6C00;
 buffer[2845] = 16'h6180;
 buffer[2846] = 16'h6023;
 buffer[2847] = 16'h710F;
 buffer[2848] = 16'h6103;
 buffer[2849] = 16'h4542;
 buffer[2850] = 16'h6E04;
 buffer[2851] = 16'h6D61;
 buffer[2852] = 16'h0065;
 buffer[2853] = 16'h0800;
 buffer[2854] = 16'h1610;
 buffer[2855] = 16'h2403;
 buffer[2856] = 16'h6E2C;
 buffer[2857] = 16'hFEBA;
 buffer[2858] = 16'h03BC;
 buffer[2859] = 16'h164E;
 buffer[2860] = 16'h2408;
 buffer[2861] = 16'h6F63;
 buffer[2862] = 16'h706D;
 buffer[2863] = 16'h6C69;
 buffer[2864] = 16'h0065;
 buffer[2865] = 16'h47A0;
 buffer[2866] = 16'h4264;
 buffer[2867] = 16'h2B3B;
 buffer[2868] = 16'h6C00;
 buffer[2869] = 16'h8080;
 buffer[2870] = 16'h6303;
 buffer[2871] = 16'h2B3A;
 buffer[2872] = 16'h0172;
 buffer[2873] = 16'h0B3B;
 buffer[2874] = 16'h08C0;
 buffer[2875] = 16'h445F;
 buffer[2876] = 16'h2B3E;
 buffer[2877] = 16'h0906;
 buffer[2878] = 16'h0800;
 buffer[2879] = 16'h1658;
 buffer[2880] = 16'h6186;
 buffer[2881] = 16'h6F62;
 buffer[2882] = 16'h7472;
 buffer[2883] = 16'h0022;
 buffer[2884] = 16'h48E6;
 buffer[2885] = 16'h480E;
 buffer[2886] = 16'h091F;
 buffer[2887] = 16'h1680;
 buffer[2888] = 16'h3C07;
 buffer[2889] = 16'h766F;
 buffer[2890] = 16'h7265;
 buffer[2891] = 16'h3E74;
 buffer[2892] = 16'hFEAE;
 buffer[2893] = 16'h6C00;
 buffer[2894] = 16'h4AE0;
 buffer[2895] = 16'h6023;
 buffer[2896] = 16'h710F;
 buffer[2897] = 16'h1690;
 buffer[2898] = 16'h6F05;
 buffer[2899] = 16'h6576;
 buffer[2900] = 16'h7472;
 buffer[2901] = 16'hFEBC;
 buffer[2902] = 16'h03BC;
 buffer[2903] = 16'h16A4;
 buffer[2904] = 16'h6504;
 buffer[2905] = 16'h6978;
 buffer[2906] = 16'h0074;
 buffer[2907] = 16'h6B8D;
 buffer[2908] = 16'h710F;
 buffer[2909] = 16'h16B0;
 buffer[2910] = 16'h3CC3;
 buffer[2911] = 16'h3E3B;
 buffer[2912] = 16'h48E6;
 buffer[2913] = 16'h4B5B;
 buffer[2914] = 16'h4847;
 buffer[2915] = 16'h4B55;
 buffer[2916] = 16'h8000;
 buffer[2917] = 16'h4394;
 buffer[2918] = 16'h6023;
 buffer[2919] = 16'h710F;
 buffer[2920] = 16'h16BC;
 buffer[2921] = 16'h3BC1;
 buffer[2922] = 16'hFEBE;
 buffer[2923] = 16'h03BC;
 buffer[2924] = 16'h16D2;
 buffer[2925] = 16'h5D01;
 buffer[2926] = 16'h9662;
 buffer[2927] = 16'hFE8A;
 buffer[2928] = 16'h6023;
 buffer[2929] = 16'h710F;
 buffer[2930] = 16'h16DA;
 buffer[2931] = 16'h3A01;
 buffer[2932] = 16'h4724;
 buffer[2933] = 16'h4B29;
 buffer[2934] = 16'h0B6E;
 buffer[2935] = 16'h16E6;
 buffer[2936] = 16'h6909;
 buffer[2937] = 16'h6D6D;
 buffer[2938] = 16'h6465;
 buffer[2939] = 16'h6169;
 buffer[2940] = 16'h6574;
 buffer[2941] = 16'h8080;
 buffer[2942] = 16'hFEAE;
 buffer[2943] = 16'h6C00;
 buffer[2944] = 16'h6C00;
 buffer[2945] = 16'h6403;
 buffer[2946] = 16'hFEAE;
 buffer[2947] = 16'h6C00;
 buffer[2948] = 16'h6023;
 buffer[2949] = 16'h710F;
 buffer[2950] = 16'h16F0;
 buffer[2951] = 16'h7504;
 buffer[2952] = 16'h6573;
 buffer[2953] = 16'h0072;
 buffer[2954] = 16'h4724;
 buffer[2955] = 16'h4B29;
 buffer[2956] = 16'h4B55;
 buffer[2957] = 16'h48E6;
 buffer[2958] = 16'h41D2;
 buffer[2959] = 16'h08B4;
 buffer[2960] = 16'h170E;
 buffer[2961] = 16'h3C08;
 buffer[2962] = 16'h7263;
 buffer[2963] = 16'h6165;
 buffer[2964] = 16'h6574;
 buffer[2965] = 16'h003E;
 buffer[2966] = 16'h4724;
 buffer[2967] = 16'h4B29;
 buffer[2968] = 16'h4B55;
 buffer[2969] = 16'h838C;
 buffer[2970] = 16'h08C0;
 buffer[2971] = 16'h1722;
 buffer[2972] = 16'h6306;
 buffer[2973] = 16'h6572;
 buffer[2974] = 16'h7461;
 buffer[2975] = 16'h0065;
 buffer[2976] = 16'hFEC0;
 buffer[2977] = 16'h03BC;
 buffer[2978] = 16'h1738;
 buffer[2979] = 16'h7608;
 buffer[2980] = 16'h7261;
 buffer[2981] = 16'h6169;
 buffer[2982] = 16'h6C62;
 buffer[2983] = 16'h0065;
 buffer[2984] = 16'h4BA0;
 buffer[2985] = 16'h8000;
 buffer[2986] = 16'h08B4;
 buffer[2987] = 16'h1746;
 buffer[2988] = 16'h3209;
 buffer[2989] = 16'h6176;
 buffer[2990] = 16'h6972;
 buffer[2991] = 16'h6261;
 buffer[2992] = 16'h656C;
 buffer[2993] = 16'h4BA0;
 buffer[2994] = 16'h8000;
 buffer[2995] = 16'h48B4;
 buffer[2996] = 16'h8001;
 buffer[2997] = 16'h4357;
 buffer[2998] = 16'h08AF;
 buffer[2999] = 16'h1758;
 buffer[3000] = 16'h2847;
 buffer[3001] = 16'h6F64;
 buffer[3002] = 16'h7365;
 buffer[3003] = 16'h293E;
 buffer[3004] = 16'h6B8D;
 buffer[3005] = 16'h8001;
 buffer[3006] = 16'h6903;
 buffer[3007] = 16'h4394;
 buffer[3008] = 16'h8001;
 buffer[3009] = 16'h6903;
 buffer[3010] = 16'hFEAE;
 buffer[3011] = 16'h6C00;
 buffer[3012] = 16'h472A;
 buffer[3013] = 16'h6081;
 buffer[3014] = 16'h434B;
 buffer[3015] = 16'hFFFF;
 buffer[3016] = 16'h6600;
 buffer[3017] = 16'h6403;
 buffer[3018] = 16'h48B4;
 buffer[3019] = 16'h6023;
 buffer[3020] = 16'h6103;
 buffer[3021] = 16'h08B4;
 buffer[3022] = 16'h1770;
 buffer[3023] = 16'h630C;
 buffer[3024] = 16'h6D6F;
 buffer[3025] = 16'h6970;
 buffer[3026] = 16'h656C;
 buffer[3027] = 16'h6F2D;
 buffer[3028] = 16'h6C6E;
 buffer[3029] = 16'h0079;
 buffer[3030] = 16'h8040;
 buffer[3031] = 16'hFEAE;
 buffer[3032] = 16'h6C00;
 buffer[3033] = 16'h6C00;
 buffer[3034] = 16'h6403;
 buffer[3035] = 16'hFEAE;
 buffer[3036] = 16'h6C00;
 buffer[3037] = 16'h6023;
 buffer[3038] = 16'h710F;
 buffer[3039] = 16'h179E;
 buffer[3040] = 16'h6485;
 buffer[3041] = 16'h656F;
 buffer[3042] = 16'h3E73;
 buffer[3043] = 16'h48E6;
 buffer[3044] = 16'h4BBC;
 buffer[3045] = 16'h700C;
 buffer[3046] = 16'h17C0;
 buffer[3047] = 16'h6304;
 buffer[3048] = 16'h6168;
 buffer[3049] = 16'h0072;
 buffer[3050] = 16'h435C;
 buffer[3051] = 16'h471C;
 buffer[3052] = 16'h6310;
 buffer[3053] = 16'h017E;
 buffer[3054] = 16'h17CE;
 buffer[3055] = 16'h5B86;
 buffer[3056] = 16'h6863;
 buffer[3057] = 16'h7261;
 buffer[3058] = 16'h005D;
 buffer[3059] = 16'h4BEA;
 buffer[3060] = 16'h0906;
 buffer[3061] = 16'h17DE;
 buffer[3062] = 16'h6308;
 buffer[3063] = 16'h6E6F;
 buffer[3064] = 16'h7473;
 buffer[3065] = 16'h6E61;
 buffer[3066] = 16'h0074;
 buffer[3067] = 16'h4BA0;
 buffer[3068] = 16'h48B4;
 buffer[3069] = 16'h4BBC;
 buffer[3070] = 16'h7C0C;
 buffer[3071] = 16'h17EC;
 buffer[3072] = 16'h6405;
 buffer[3073] = 16'h6665;
 buffer[3074] = 16'h7265;
 buffer[3075] = 16'h4BA0;
 buffer[3076] = 16'h8000;
 buffer[3077] = 16'h48B4;
 buffer[3078] = 16'h4BBC;
 buffer[3079] = 16'h6C00;
 buffer[3080] = 16'h4264;
 buffer[3081] = 16'h8000;
 buffer[3082] = 16'h6703;
 buffer[3083] = 16'h480E;
 buffer[3084] = 16'h750D;
 buffer[3085] = 16'h696E;
 buffer[3086] = 16'h696E;
 buffer[3087] = 16'h6974;
 buffer[3088] = 16'h6C61;
 buffer[3089] = 16'h7A69;
 buffer[3090] = 16'h6465;
 buffer[3091] = 16'h0172;
 buffer[3092] = 16'h1800;
 buffer[3093] = 16'h6982;
 buffer[3094] = 16'h0073;
 buffer[3095] = 16'h48A6;
 buffer[3096] = 16'h4AB3;
 buffer[3097] = 16'h6023;
 buffer[3098] = 16'h710F;
 buffer[3099] = 16'h182A;
 buffer[3100] = 16'h2E03;
 buffer[3101] = 16'h6469;
 buffer[3102] = 16'h4264;
 buffer[3103] = 16'h2C24;
 buffer[3104] = 16'h438C;
 buffer[3105] = 16'h801F;
 buffer[3106] = 16'h6303;
 buffer[3107] = 16'h051E;
 buffer[3108] = 16'h452E;
 buffer[3109] = 16'h454C;
 buffer[3110] = 16'h7B08;
 buffer[3111] = 16'h6F6E;
 buffer[3112] = 16'h616E;
 buffer[3113] = 16'h656D;
 buffer[3114] = 16'h007D;
 buffer[3115] = 16'h700C;
 buffer[3116] = 16'h1838;
 buffer[3117] = 16'h7708;
 buffer[3118] = 16'h726F;
 buffer[3119] = 16'h6C64;
 buffer[3120] = 16'h7369;
 buffer[3121] = 16'h0074;
 buffer[3122] = 16'h43AA;
 buffer[3123] = 16'h4394;
 buffer[3124] = 16'h8000;
 buffer[3125] = 16'h48B4;
 buffer[3126] = 16'h6081;
 buffer[3127] = 16'hFEA8;
 buffer[3128] = 16'h434B;
 buffer[3129] = 16'h6081;
 buffer[3130] = 16'h6C00;
 buffer[3131] = 16'h48B4;
 buffer[3132] = 16'h6023;
 buffer[3133] = 16'h6103;
 buffer[3134] = 16'h8000;
 buffer[3135] = 16'h08B4;
 buffer[3136] = 16'h185A;
 buffer[3137] = 16'h6F06;
 buffer[3138] = 16'h6472;
 buffer[3139] = 16'h7265;
 buffer[3140] = 16'h0040;
 buffer[3141] = 16'h6081;
 buffer[3142] = 16'h6C00;
 buffer[3143] = 16'h6081;
 buffer[3144] = 16'h2C4F;
 buffer[3145] = 16'h6147;
 buffer[3146] = 16'h434B;
 buffer[3147] = 16'h4C45;
 buffer[3148] = 16'h6B8D;
 buffer[3149] = 16'h6180;
 buffer[3150] = 16'h731C;
 buffer[3151] = 16'h700F;
 buffer[3152] = 16'h1882;
 buffer[3153] = 16'h6709;
 buffer[3154] = 16'h7465;
 buffer[3155] = 16'h6F2D;
 buffer[3156] = 16'h6472;
 buffer[3157] = 16'h7265;
 buffer[3158] = 16'hFE90;
 buffer[3159] = 16'h0C45;
 buffer[3160] = 16'h18A2;
 buffer[3161] = 16'h3E04;
 buffer[3162] = 16'h6977;
 buffer[3163] = 16'h0064;
 buffer[3164] = 16'h034B;
 buffer[3165] = 16'h18B2;
 buffer[3166] = 16'h2E04;
 buffer[3167] = 16'h6977;
 buffer[3168] = 16'h0064;
 buffer[3169] = 16'h4506;
 buffer[3170] = 16'h6081;
 buffer[3171] = 16'h4C5C;
 buffer[3172] = 16'h434B;
 buffer[3173] = 16'h6C00;
 buffer[3174] = 16'h4264;
 buffer[3175] = 16'h2C6A;
 buffer[3176] = 16'h4C1E;
 buffer[3177] = 16'h710F;
 buffer[3178] = 16'h8000;
 buffer[3179] = 16'h055B;
 buffer[3180] = 16'h18BC;
 buffer[3181] = 16'h2104;
 buffer[3182] = 16'h6977;
 buffer[3183] = 16'h0064;
 buffer[3184] = 16'h4C5C;
 buffer[3185] = 16'h434B;
 buffer[3186] = 16'hFEAE;
 buffer[3187] = 16'h6C00;
 buffer[3188] = 16'h6180;
 buffer[3189] = 16'h6023;
 buffer[3190] = 16'h710F;
 buffer[3191] = 16'h18DA;
 buffer[3192] = 16'h7604;
 buffer[3193] = 16'h636F;
 buffer[3194] = 16'h0073;
 buffer[3195] = 16'h452E;
 buffer[3196] = 16'h454C;
 buffer[3197] = 16'h7605;
 buffer[3198] = 16'h636F;
 buffer[3199] = 16'h3A73;
 buffer[3200] = 16'hFEA8;
 buffer[3201] = 16'h434B;
 buffer[3202] = 16'h6C00;
 buffer[3203] = 16'h4264;
 buffer[3204] = 16'h2C89;
 buffer[3205] = 16'h6081;
 buffer[3206] = 16'h4C61;
 buffer[3207] = 16'h4C5C;
 buffer[3208] = 16'h0C82;
 buffer[3209] = 16'h700C;
 buffer[3210] = 16'h18F0;
 buffer[3211] = 16'h6F05;
 buffer[3212] = 16'h6472;
 buffer[3213] = 16'h7265;
 buffer[3214] = 16'h452E;
 buffer[3215] = 16'h454C;
 buffer[3216] = 16'h7307;
 buffer[3217] = 16'h6165;
 buffer[3218] = 16'h6372;
 buffer[3219] = 16'h3A68;
 buffer[3220] = 16'h4C56;
 buffer[3221] = 16'h4264;
 buffer[3222] = 16'h2C9B;
 buffer[3223] = 16'h6180;
 buffer[3224] = 16'h4C61;
 buffer[3225] = 16'h6A00;
 buffer[3226] = 16'h0C95;
 buffer[3227] = 16'h452E;
 buffer[3228] = 16'h454C;
 buffer[3229] = 16'h6407;
 buffer[3230] = 16'h6665;
 buffer[3231] = 16'h6E69;
 buffer[3232] = 16'h3A65;
 buffer[3233] = 16'h4AE0;
 buffer[3234] = 16'h0C61;
 buffer[3235] = 16'h1916;
 buffer[3236] = 16'h7309;
 buffer[3237] = 16'h7465;
 buffer[3238] = 16'h6F2D;
 buffer[3239] = 16'h6472;
 buffer[3240] = 16'h7265;
 buffer[3241] = 16'h6081;
 buffer[3242] = 16'h8000;
 buffer[3243] = 16'h6600;
 buffer[3244] = 16'h6703;
 buffer[3245] = 16'h2CB1;
 buffer[3246] = 16'h6103;
 buffer[3247] = 16'hFEA2;
 buffer[3248] = 16'h8001;
 buffer[3249] = 16'h8008;
 buffer[3250] = 16'h6181;
 buffer[3251] = 16'h6F03;
 buffer[3252] = 16'h480E;
 buffer[3253] = 16'h6F12;
 buffer[3254] = 16'h6576;
 buffer[3255] = 16'h2072;
 buffer[3256] = 16'h6973;
 buffer[3257] = 16'h657A;
 buffer[3258] = 16'h6F20;
 buffer[3259] = 16'h2066;
 buffer[3260] = 16'h7623;
 buffer[3261] = 16'h636F;
 buffer[3262] = 16'h0073;
 buffer[3263] = 16'hFE90;
 buffer[3264] = 16'h6180;
 buffer[3265] = 16'h6081;
 buffer[3266] = 16'h2CCC;
 buffer[3267] = 16'h6147;
 buffer[3268] = 16'h6180;
 buffer[3269] = 16'h6181;
 buffer[3270] = 16'h6023;
 buffer[3271] = 16'h6103;
 buffer[3272] = 16'h434B;
 buffer[3273] = 16'h6B8D;
 buffer[3274] = 16'h6A00;
 buffer[3275] = 16'h0CC1;
 buffer[3276] = 16'h6180;
 buffer[3277] = 16'h6023;
 buffer[3278] = 16'h710F;
 buffer[3279] = 16'h1948;
 buffer[3280] = 16'h6F04;
 buffer[3281] = 16'h6C6E;
 buffer[3282] = 16'h0079;
 buffer[3283] = 16'h8000;
 buffer[3284] = 16'h6600;
 buffer[3285] = 16'h0CA9;
 buffer[3286] = 16'h19A0;
 buffer[3287] = 16'h6104;
 buffer[3288] = 16'h736C;
 buffer[3289] = 16'h006F;
 buffer[3290] = 16'h4C56;
 buffer[3291] = 16'h6181;
 buffer[3292] = 16'h6180;
 buffer[3293] = 16'h6310;
 buffer[3294] = 16'h0CA9;
 buffer[3295] = 16'h19AE;
 buffer[3296] = 16'h7008;
 buffer[3297] = 16'h6572;
 buffer[3298] = 16'h6976;
 buffer[3299] = 16'h756F;
 buffer[3300] = 16'h0073;
 buffer[3301] = 16'h4C56;
 buffer[3302] = 16'h6180;
 buffer[3303] = 16'h6103;
 buffer[3304] = 16'h6A00;
 buffer[3305] = 16'h0CA9;
 buffer[3306] = 16'h19C0;
 buffer[3307] = 16'h3E04;
 buffer[3308] = 16'h6F76;
 buffer[3309] = 16'h0063;
 buffer[3310] = 16'h4BA0;
 buffer[3311] = 16'h6081;
 buffer[3312] = 16'h48B4;
 buffer[3313] = 16'h4C70;
 buffer[3314] = 16'h4BBC;
 buffer[3315] = 16'h6C00;
 buffer[3316] = 16'h6147;
 buffer[3317] = 16'h4C56;
 buffer[3318] = 16'h6180;
 buffer[3319] = 16'h6103;
 buffer[3320] = 16'h6B8D;
 buffer[3321] = 16'h6180;
 buffer[3322] = 16'h0CA9;
 buffer[3323] = 16'h19D6;
 buffer[3324] = 16'h7705;
 buffer[3325] = 16'h6469;
 buffer[3326] = 16'h666F;
 buffer[3327] = 16'h48A6;
 buffer[3328] = 16'h4AB3;
 buffer[3329] = 16'h7C0C;
 buffer[3330] = 16'h19F8;
 buffer[3331] = 16'h760A;
 buffer[3332] = 16'h636F;
 buffer[3333] = 16'h6261;
 buffer[3334] = 16'h6C75;
 buffer[3335] = 16'h7261;
 buffer[3336] = 16'h0079;
 buffer[3337] = 16'h4C32;
 buffer[3338] = 16'h0CEE;
 buffer[3339] = 16'h1A06;
 buffer[3340] = 16'h5F05;
 buffer[3341] = 16'h7974;
 buffer[3342] = 16'h6570;
 buffer[3343] = 16'h6147;
 buffer[3344] = 16'h0D14;
 buffer[3345] = 16'h438C;
 buffer[3346] = 16'h4362;
 buffer[3347] = 16'h44CC;
 buffer[3348] = 16'h6B81;
 buffer[3349] = 16'h2D1A;
 buffer[3350] = 16'h6B8D;
 buffer[3351] = 16'h6A00;
 buffer[3352] = 16'h6147;
 buffer[3353] = 16'h0D11;
 buffer[3354] = 16'h6B8D;
 buffer[3355] = 16'h6103;
 buffer[3356] = 16'h710F;
 buffer[3357] = 16'h1A18;
 buffer[3358] = 16'h6403;
 buffer[3359] = 16'h2B6D;
 buffer[3360] = 16'h6181;
 buffer[3361] = 16'h8004;
 buffer[3362] = 16'h455B;
 buffer[3363] = 16'h4506;
 buffer[3364] = 16'h6147;
 buffer[3365] = 16'h0D29;
 buffer[3366] = 16'h438C;
 buffer[3367] = 16'h8003;
 buffer[3368] = 16'h455B;
 buffer[3369] = 16'h6B81;
 buffer[3370] = 16'h2D2F;
 buffer[3371] = 16'h6B8D;
 buffer[3372] = 16'h6A00;
 buffer[3373] = 16'h6147;
 buffer[3374] = 16'h0D26;
 buffer[3375] = 16'h6B8D;
 buffer[3376] = 16'h710F;
 buffer[3377] = 16'h1A3C;
 buffer[3378] = 16'h6404;
 buffer[3379] = 16'h6D75;
 buffer[3380] = 16'h0070;
 buffer[3381] = 16'hFE80;
 buffer[3382] = 16'h6C00;
 buffer[3383] = 16'h6147;
 buffer[3384] = 16'h4432;
 buffer[3385] = 16'h8010;
 buffer[3386] = 16'h4305;
 buffer[3387] = 16'h6147;
 buffer[3388] = 16'h452E;
 buffer[3389] = 16'h8010;
 buffer[3390] = 16'h4279;
 buffer[3391] = 16'h4D20;
 buffer[3392] = 16'h4155;
 buffer[3393] = 16'h8002;
 buffer[3394] = 16'h450D;
 buffer[3395] = 16'h4D0F;
 buffer[3396] = 16'h6B81;
 buffer[3397] = 16'h2D4A;
 buffer[3398] = 16'h6B8D;
 buffer[3399] = 16'h6A00;
 buffer[3400] = 16'h6147;
 buffer[3401] = 16'h0D3C;
 buffer[3402] = 16'h6B8D;
 buffer[3403] = 16'h6103;
 buffer[3404] = 16'h6103;
 buffer[3405] = 16'h6B8D;
 buffer[3406] = 16'hFE80;
 buffer[3407] = 16'h6023;
 buffer[3408] = 16'h710F;
 buffer[3409] = 16'h1A64;
 buffer[3410] = 16'h2E02;
 buffer[3411] = 16'h0073;
 buffer[3412] = 16'h452E;
 buffer[3413] = 16'h416A;
 buffer[3414] = 16'h6A00;
 buffer[3415] = 16'h800F;
 buffer[3416] = 16'h6303;
 buffer[3417] = 16'h6147;
 buffer[3418] = 16'h6B81;
 buffer[3419] = 16'h48FA;
 buffer[3420] = 16'h456E;
 buffer[3421] = 16'h6B81;
 buffer[3422] = 16'h2D63;
 buffer[3423] = 16'h6B8D;
 buffer[3424] = 16'h6A00;
 buffer[3425] = 16'h6147;
 buffer[3426] = 16'h0D5A;
 buffer[3427] = 16'h6B8D;
 buffer[3428] = 16'h6103;
 buffer[3429] = 16'h454C;
 buffer[3430] = 16'h3C04;
 buffer[3431] = 16'h6F74;
 buffer[3432] = 16'h0073;
 buffer[3433] = 16'h700C;
 buffer[3434] = 16'h1AA4;
 buffer[3435] = 16'h2807;
 buffer[3436] = 16'h6E3E;
 buffer[3437] = 16'h6D61;
 buffer[3438] = 16'h2965;
 buffer[3439] = 16'h6C00;
 buffer[3440] = 16'h4264;
 buffer[3441] = 16'h2D79;
 buffer[3442] = 16'h4279;
 buffer[3443] = 16'h472A;
 buffer[3444] = 16'h6503;
 buffer[3445] = 16'h2D78;
 buffer[3446] = 16'h4351;
 buffer[3447] = 16'h0D6F;
 buffer[3448] = 16'h700F;
 buffer[3449] = 16'h6103;
 buffer[3450] = 16'h8000;
 buffer[3451] = 16'h700C;
 buffer[3452] = 16'h1AD6;
 buffer[3453] = 16'h3E05;
 buffer[3454] = 16'h616E;
 buffer[3455] = 16'h656D;
 buffer[3456] = 16'h6147;
 buffer[3457] = 16'h4C56;
 buffer[3458] = 16'h4264;
 buffer[3459] = 16'h2D9C;
 buffer[3460] = 16'h6180;
 buffer[3461] = 16'h6B81;
 buffer[3462] = 16'h6180;
 buffer[3463] = 16'h4D6F;
 buffer[3464] = 16'h4264;
 buffer[3465] = 16'h2D9A;
 buffer[3466] = 16'h6147;
 buffer[3467] = 16'h6A00;
 buffer[3468] = 16'h6147;
 buffer[3469] = 16'h0D8F;
 buffer[3470] = 16'h6103;
 buffer[3471] = 16'h6B81;
 buffer[3472] = 16'h2D95;
 buffer[3473] = 16'h6B8D;
 buffer[3474] = 16'h6A00;
 buffer[3475] = 16'h6147;
 buffer[3476] = 16'h0D8E;
 buffer[3477] = 16'h6B8D;
 buffer[3478] = 16'h6103;
 buffer[3479] = 16'h6B8D;
 buffer[3480] = 16'h6B8D;
 buffer[3481] = 16'h710F;
 buffer[3482] = 16'h6A00;
 buffer[3483] = 16'h0D82;
 buffer[3484] = 16'h6B8D;
 buffer[3485] = 16'h6103;
 buffer[3486] = 16'h8000;
 buffer[3487] = 16'h700C;
 buffer[3488] = 16'h1AFA;
 buffer[3489] = 16'h7303;
 buffer[3490] = 16'h6565;
 buffer[3491] = 16'h48A6;
 buffer[3492] = 16'h452E;
 buffer[3493] = 16'h6081;
 buffer[3494] = 16'h6C00;
 buffer[3495] = 16'h4264;
 buffer[3496] = 16'hF00C;
 buffer[3497] = 16'h6503;
 buffer[3498] = 16'h2DBC;
 buffer[3499] = 16'hBFFF;
 buffer[3500] = 16'h6303;
 buffer[3501] = 16'h8001;
 buffer[3502] = 16'h6D03;
 buffer[3503] = 16'h4D80;
 buffer[3504] = 16'h4264;
 buffer[3505] = 16'h2DB5;
 buffer[3506] = 16'h4506;
 buffer[3507] = 16'h4C1E;
 buffer[3508] = 16'h0DBA;
 buffer[3509] = 16'h6081;
 buffer[3510] = 16'h6C00;
 buffer[3511] = 16'hFFFF;
 buffer[3512] = 16'h6303;
 buffer[3513] = 16'h4567;
 buffer[3514] = 16'h434B;
 buffer[3515] = 16'h0DA5;
 buffer[3516] = 16'h0273;
 buffer[3517] = 16'h1B42;
 buffer[3518] = 16'h2807;
 buffer[3519] = 16'h6F77;
 buffer[3520] = 16'h6472;
 buffer[3521] = 16'h2973;
 buffer[3522] = 16'h452E;
 buffer[3523] = 16'h6C00;
 buffer[3524] = 16'h4264;
 buffer[3525] = 16'h2DCB;
 buffer[3526] = 16'h6081;
 buffer[3527] = 16'h4C1E;
 buffer[3528] = 16'h4506;
 buffer[3529] = 16'h4351;
 buffer[3530] = 16'h0DC3;
 buffer[3531] = 16'h700C;
 buffer[3532] = 16'h1B7C;
 buffer[3533] = 16'h7705;
 buffer[3534] = 16'h726F;
 buffer[3535] = 16'h7364;
 buffer[3536] = 16'h4C56;
 buffer[3537] = 16'h4264;
 buffer[3538] = 16'h2DDE;
 buffer[3539] = 16'h6180;
 buffer[3540] = 16'h452E;
 buffer[3541] = 16'h452E;
 buffer[3542] = 16'h454C;
 buffer[3543] = 16'h3A01;
 buffer[3544] = 16'h6081;
 buffer[3545] = 16'h4C61;
 buffer[3546] = 16'h452E;
 buffer[3547] = 16'h4DC2;
 buffer[3548] = 16'h6A00;
 buffer[3549] = 16'h0DD1;
 buffer[3550] = 16'h700C;
 buffer[3551] = 16'h1B9A;
 buffer[3552] = 16'h7603;
 buffer[3553] = 16'h7265;
 buffer[3554] = 16'h8001;
 buffer[3555] = 16'h8100;
 buffer[3556] = 16'h4329;
 buffer[3557] = 16'h8006;
 buffer[3558] = 16'h720F;
 buffer[3559] = 16'h1BC0;
 buffer[3560] = 16'h6802;
 buffer[3561] = 16'h0069;
 buffer[3562] = 16'h452E;
 buffer[3563] = 16'h454C;
 buffer[3564] = 16'h650C;
 buffer[3565] = 16'h6F66;
 buffer[3566] = 16'h7472;
 buffer[3567] = 16'h2068;
 buffer[3568] = 16'h316A;
 buffer[3569] = 16'h202B;
 buffer[3570] = 16'h0076;
 buffer[3571] = 16'hFE80;
 buffer[3572] = 16'h6C00;
 buffer[3573] = 16'h4432;
 buffer[3574] = 16'h4DE2;
 buffer[3575] = 16'h43F4;
 buffer[3576] = 16'h4406;
 buffer[3577] = 16'h4406;
 buffer[3578] = 16'h802E;
 buffer[3579] = 16'h43FC;
 buffer[3580] = 16'h4406;
 buffer[3581] = 16'h441E;
 buffer[3582] = 16'h451E;
 buffer[3583] = 16'hFE80;
 buffer[3584] = 16'h6023;
 buffer[3585] = 16'h6103;
 buffer[3586] = 16'h052E;
 buffer[3587] = 16'h1BD0;
 buffer[3588] = 16'h6304;
 buffer[3589] = 16'h6C6F;
 buffer[3590] = 16'h0064;
 buffer[3591] = 16'h8002;
 buffer[3592] = 16'hFE80;
 buffer[3593] = 16'h8042;
 buffer[3594] = 16'h45BC;
 buffer[3595] = 16'h488E;
 buffer[3596] = 16'hFEA2;
 buffer[3597] = 16'h6081;
 buffer[3598] = 16'hFE90;
 buffer[3599] = 16'h6023;
 buffer[3600] = 16'h6103;
 buffer[3601] = 16'h6081;
 buffer[3602] = 16'hFEA8;
 buffer[3603] = 16'h4379;
 buffer[3604] = 16'h4B55;
 buffer[3605] = 16'hC000;
 buffer[3606] = 16'h434B;
 buffer[3607] = 16'h6081;
 buffer[3608] = 16'h4351;
 buffer[3609] = 16'h6C00;
 buffer[3610] = 16'h4868;
 buffer[3611] = 16'hFEB4;
 buffer[3612] = 16'h43BC;
 buffer[3613] = 16'h4897;
 buffer[3614] = 16'h0E07;
end

endmodule

module M_main_mem_ram(
input      [0:0]             in_ram_wenable0,
input       [15:0]     in_ram_wdata0,
input      [14:0]                in_ram_addr0,
input      [0:0]             in_ram_wenable1,
input      [15:0]                 in_ram_wdata1,
input      [14:0]                in_ram_addr1,
output reg  [15:0]     out_ram_rdata0,
output reg  [15:0]     out_ram_rdata1,
input      clock0,
input      clock1
);
reg  [15:0] buffer[32767:0];
always @(posedge clock0) begin
  if (in_ram_wenable0) begin
    buffer[in_ram_addr0] <= in_ram_wdata0;
  end else begin
    out_ram_rdata0 <= buffer[in_ram_addr0];
  end
end
always @(posedge clock1) begin
  if (in_ram_wenable1) begin
    buffer[in_ram_addr1] <= in_ram_wdata1;
  end else begin
    out_ram_rdata1 <= buffer[in_ram_addr1];
  end
end

endmodule

module M_main_mem_uartInBuffer(
input      [0:0]             in_uartInBuffer_wenable0,
input       [7:0]     in_uartInBuffer_wdata0,
input      [8:0]                in_uartInBuffer_addr0,
input      [0:0]             in_uartInBuffer_wenable1,
input      [7:0]                 in_uartInBuffer_wdata1,
input      [8:0]                in_uartInBuffer_addr1,
output reg  [7:0]     out_uartInBuffer_rdata0,
output reg  [7:0]     out_uartInBuffer_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[511:0];
always @(posedge clock0) begin
  if (in_uartInBuffer_wenable0) begin
    buffer[in_uartInBuffer_addr0] <= in_uartInBuffer_wdata0;
  end else begin
    out_uartInBuffer_rdata0 <= buffer[in_uartInBuffer_addr0];
  end
end
always @(posedge clock1) begin
  if (in_uartInBuffer_wenable1) begin
    buffer[in_uartInBuffer_addr1] <= in_uartInBuffer_wdata1;
  end else begin
    out_uartInBuffer_rdata1 <= buffer[in_uartInBuffer_addr1];
  end
end

endmodule

module M_main_mem_uartOutBuffer(
input      [0:0]             in_uartOutBuffer_wenable0,
input       [7:0]     in_uartOutBuffer_wdata0,
input      [8:0]                in_uartOutBuffer_addr0,
input      [0:0]             in_uartOutBuffer_wenable1,
input      [7:0]                 in_uartOutBuffer_wdata1,
input      [8:0]                in_uartOutBuffer_addr1,
output reg  [7:0]     out_uartOutBuffer_rdata0,
output reg  [7:0]     out_uartOutBuffer_rdata1,
input      clock0,
input      clock1
);
reg  [7:0] buffer[511:0];
always @(posedge clock0) begin
  if (in_uartOutBuffer_wenable0) begin
    buffer[in_uartOutBuffer_addr0] <= in_uartOutBuffer_wdata0;
  end else begin
    out_uartOutBuffer_rdata0 <= buffer[in_uartOutBuffer_addr0];
  end
end
always @(posedge clock1) begin
  if (in_uartOutBuffer_wenable1) begin
    buffer[in_uartOutBuffer_addr1] <= in_uartOutBuffer_wdata1;
  end else begin
    out_uartOutBuffer_rdata1 <= buffer[in_uartOutBuffer_addr1];
  end
end

endmodule

module M_main (
in_buttons,
in_uart_tx_busy,
in_uart_tx_done,
in_uart_rx_data,
in_uart_rx_valid,
in_timer1hz,
out_led,
out_uart_tx_data,
out_uart_tx_valid,
out_uart_rx_ready,
out_sdram_cle,
out_sdram_dqm,
out_sdram_cs,
out_sdram_we,
out_sdram_cas,
out_sdram_ras,
out_sdram_ba,
out_sdram_a,
out_sdram_clk,
out_video_r,
out_video_g,
out_video_b,
out_video_hs,
out_video_vs,
inout_sdram_dq,
in_run,
out_done,
reset,
clock
);
input  [7:0] in_buttons;
input  [0:0] in_uart_tx_busy;
input  [0:0] in_uart_tx_done;
input  [7:0] in_uart_rx_data;
input  [0:0] in_uart_rx_valid;
input  [15:0] in_timer1hz;
output  [7:0] out_led;
output  [7:0] out_uart_tx_data;
output  [0:0] out_uart_tx_valid;
output  [0:0] out_uart_rx_ready;
output  [0:0] out_sdram_cle;
output  [0:0] out_sdram_dqm;
output  [0:0] out_sdram_cs;
output  [0:0] out_sdram_we;
output  [0:0] out_sdram_cas;
output  [0:0] out_sdram_ras;
output  [1:0] out_sdram_ba;
output  [12:0] out_sdram_a;
output  [0:0] out_sdram_clk;
output  [5:0] out_video_r;
output  [5:0] out_video_g;
output  [5:0] out_video_b;
output  [0:0] out_video_hs;
output  [0:0] out_video_vs;
inout  [7:0] inout_sdram_dq;
input in_run;
output out_done;
input reset;
input clock;
wire _w_vga_rstcond_out;
wire _w_clk_gen_outclk_0;
wire _w_clk_gen_outclk_1;
wire _w_clk_gen_locked;
wire  [0:0] _w_vga_driver_vga_hs;
wire  [0:0] _w_vga_driver_vga_vs;
wire  [0:0] _w_vga_driver_active;
wire  [0:0] _w_vga_driver_vblank;
wire  [9:0] _w_vga_driver_vga_x;
wire  [9:0] _w_vga_driver_vga_y;
wire _w_vga_driver_done;
wire  [5:0] _w_display_pix_red;
wire  [5:0] _w_display_pix_green;
wire  [5:0] _w_display_pix_blue;
wire  [7:0] _w_display_gpu_active;
wire _w_display_done;
wire  [15:0] _w_mem_dstack_rdata;
wire  [15:0] _w_mem_rstack_rdata;
wire  [15:0] _w_mem_rom_rdata;
wire  [15:0] _w_mem_ram_rdata0;
wire  [15:0] _w_mem_ram_rdata1;
wire  [7:0] _w_mem_uartInBuffer_rdata0;
wire  [7:0] _w_mem_uartInBuffer_rdata1;
wire  [7:0] _w_mem_uartOutBuffer_rdata0;
wire  [7:0] _w_mem_uartOutBuffer_rdata1;
wire  [15:0] _c_ram_wdata1;
assign _c_ram_wdata1 = 0;
wire  [7:0] _c_uartInBuffer_wdata0;
assign _c_uartInBuffer_wdata0 = 0;
wire  [7:0] _c_uartOutBuffer_wdata0;
assign _c_uartOutBuffer_wdata0 = 0;
wire  [15:0] _w_immediate;
wire  [0:0] _w_is_alu;
wire  [0:0] _w_is_call;
wire  [0:0] _w_is_lit;
wire  [0:0] _w_dstackWrite;
wire  [0:0] _w_rstackWrite;
wire  [7:0] _w_ddelta;
wire  [7:0] _w_rdelta;
wire  [12:0] _w_pcPlusOne;

reg  [15:0] _d_instruction;
reg  [15:0] _q_instruction;
reg  [12:0] _d_pc;
reg  [12:0] _q_pc;
reg  [12:0] _d_newPC;
reg  [12:0] _q_newPC;
reg  [0:0] _d_dstack_wenable;
reg  [0:0] _q_dstack_wenable;
reg  [15:0] _d_dstack_wdata;
reg  [15:0] _q_dstack_wdata;
reg  [7:0] _d_dstack_addr;
reg  [7:0] _q_dstack_addr;
reg  [15:0] _d_stackTop;
reg  [15:0] _q_stackTop;
reg  [7:0] _d_dsp;
reg  [7:0] _q_dsp;
reg  [7:0] _d_newDSP;
reg  [7:0] _q_newDSP;
reg  [15:0] _d_newStackTop;
reg  [15:0] _q_newStackTop;
reg  [0:0] _d_rstack_wenable;
reg  [0:0] _q_rstack_wenable;
reg  [15:0] _d_rstack_wdata;
reg  [15:0] _q_rstack_wdata;
reg  [7:0] _d_rstack_addr;
reg  [7:0] _q_rstack_addr;
reg  [7:0] _d_rsp;
reg  [7:0] _q_rsp;
reg  [7:0] _d_newRSP;
reg  [7:0] _q_newRSP;
reg  [15:0] _d_rstackWData;
reg  [15:0] _q_rstackWData;
reg  [15:0] _d_stackNext;
reg  [15:0] _q_stackNext;
reg  [15:0] _d_rStackTop;
reg  [15:0] _q_rStackTop;
reg  [15:0] _d_memoryInput;
reg  [15:0] _q_memoryInput;
reg  [11:0] _d_rom_addr;
reg  [11:0] _q_rom_addr;
reg  [0:0] _d_ram_wenable0;
reg  [0:0] _q_ram_wenable0;
reg  [15:0] _d_ram_wdata0;
reg  [15:0] _q_ram_wdata0;
reg  [14:0] _d_ram_addr0;
reg  [14:0] _q_ram_addr0;
reg  [0:0] _d_ram_wenable1;
reg  [0:0] _q_ram_wenable1;
reg  [14:0] _d_ram_addr1;
reg  [14:0] _q_ram_addr1;
reg  [2:0] _d_CYCLE;
reg  [2:0] _q_CYCLE;
reg  [1:0] _d_INIT;
reg  [1:0] _q_INIT;
reg  [15:0] _d_copyaddress;
reg  [15:0] _q_copyaddress;
reg  [15:0] _d_bramREAD;
reg  [15:0] _q_bramREAD;
reg  [0:0] _d_uartInBuffer_wenable0;
reg  [0:0] _q_uartInBuffer_wenable0;
reg  [8:0] _d_uartInBuffer_addr0;
reg  [8:0] _q_uartInBuffer_addr0;
reg  [0:0] _d_uartInBuffer_wenable1;
reg  [0:0] _q_uartInBuffer_wenable1;
reg  [7:0] _d_uartInBuffer_wdata1;
reg  [7:0] _q_uartInBuffer_wdata1;
reg  [8:0] _d_uartInBuffer_addr1;
reg  [8:0] _q_uartInBuffer_addr1;
reg  [8:0] _d_uartInBufferNext;
reg  [8:0] _q_uartInBufferNext;
reg  [8:0] _d_uartInBufferTop;
reg  [8:0] _q_uartInBufferTop;
reg  [0:0] _d_uartInHold;
reg  [0:0] _q_uartInHold;
reg  [0:0] _d_uartOutBuffer_wenable0;
reg  [0:0] _q_uartOutBuffer_wenable0;
reg  [8:0] _d_uartOutBuffer_addr0;
reg  [8:0] _q_uartOutBuffer_addr0;
reg  [0:0] _d_uartOutBuffer_wenable1;
reg  [0:0] _q_uartOutBuffer_wenable1;
reg  [7:0] _d_uartOutBuffer_wdata1;
reg  [7:0] _q_uartOutBuffer_wdata1;
reg  [8:0] _d_uartOutBuffer_addr1;
reg  [8:0] _q_uartOutBuffer_addr1;
reg  [8:0] _d_uartOutBufferNext;
reg  [8:0] _q_uartOutBufferNext;
reg  [8:0] _d_uartOutBufferTop;
reg  [8:0] _q_uartOutBufferTop;
reg  [8:0] _d_newuartOutBufferTop;
reg  [8:0] _q_newuartOutBufferTop;
reg  [0:0] _d_uartOutHold;
reg  [0:0] _q_uartOutHold;
reg  [7:0] _d_led,_q_led;
reg  [7:0] _d_uart_tx_data,_q_uart_tx_data;
reg  [0:0] _d_uart_tx_valid,_q_uart_tx_valid;
reg  [0:0] _d_uart_rx_ready,_q_uart_rx_ready;
reg  [0:0] _d_sdram_cle,_q_sdram_cle;
reg  [0:0] _d_sdram_dqm,_q_sdram_dqm;
reg  [0:0] _d_sdram_cs,_q_sdram_cs;
reg  [0:0] _d_sdram_we,_q_sdram_we;
reg  [0:0] _d_sdram_cas,_q_sdram_cas;
reg  [0:0] _d_sdram_ras,_q_sdram_ras;
reg  [1:0] _d_sdram_ba,_q_sdram_ba;
reg  [12:0] _d_sdram_a,_q_sdram_a;
reg  [0:0] _d_sdram_clk,_q_sdram_clk;
reg  [9:0] _d_display_gpu_x,_q_display_gpu_x;
reg  [8:0] _d_display_gpu_y,_q_display_gpu_y;
reg  [15:0] _d_display_gpu_param0,_q_display_gpu_param0;
reg  [15:0] _d_display_gpu_param1,_q_display_gpu_param1;
reg  [15:0] _d_display_gpu_param2,_q_display_gpu_param2;
reg  [15:0] _d_display_gpu_param3,_q_display_gpu_param3;
reg  [7:0] _d_display_gpu_colour,_q_display_gpu_colour;
reg  [1:0] _d_display_gpu_write,_q_display_gpu_write;
reg  [6:0] _d_display_tpu_x,_q_display_tpu_x;
reg  [4:0] _d_display_tpu_y,_q_display_tpu_y;
reg  [7:0] _d_display_tpu_set,_q_display_tpu_set;
reg  [1:0] _d_display_tpu_write,_q_display_tpu_write;
reg  [7:0] _d_display_terminal_character,_q_display_terminal_character;
reg  [0:0] _d_display_terminal_write,_q_display_terminal_write;
reg  [0:0] _d_display_showterminal,_q_display_showterminal;
reg  [0:0] _d_display_showcursor,_q_display_showcursor;
reg  [2:0] _d_index,_q_index;
reg  _vga_driver_run;
reg  _display_run;
assign out_led = _q_led;
assign out_uart_tx_data = _q_uart_tx_data;
assign out_uart_tx_valid = _q_uart_tx_valid;
assign out_uart_rx_ready = _q_uart_rx_ready;
assign out_sdram_cle = _d_sdram_cle;
assign out_sdram_dqm = _d_sdram_dqm;
assign out_sdram_cs = _d_sdram_cs;
assign out_sdram_we = _d_sdram_we;
assign out_sdram_cas = _d_sdram_cas;
assign out_sdram_ras = _d_sdram_ras;
assign out_sdram_ba = _d_sdram_ba;
assign out_sdram_a = _d_sdram_a;
assign out_sdram_clk = _d_sdram_clk;
assign out_video_r = _w_display_pix_red;
assign out_video_g = _w_display_pix_green;
assign out_video_b = _w_display_pix_blue;
assign out_video_hs = _w_vga_driver_vga_hs;
assign out_video_vs = _w_vga_driver_vga_vs;
assign out_done = (_q_index == 7);

always @(posedge clock) begin
  if (reset || !in_run) begin
_q_pc <= 0;
_q_dstack_wenable <= 0;
_q_dstack_wdata <= 0;
_q_dstack_addr <= 0;
_q_stackTop <= 0;
_q_dsp <= 0;
_q_rstack_wenable <= 0;
_q_rstack_wdata <= 0;
_q_rstack_addr <= 0;
_q_rsp <= 0;
_q_rom_addr <= 0;
_q_ram_wenable0 <= 0;
_q_ram_wdata0 <= 0;
_q_ram_addr0 <= 0;
_q_ram_wenable1 <= 0;
_q_ram_addr1 <= 0;
_q_CYCLE <= 0;
_q_INIT <= 0;
_q_copyaddress <= 0;
_q_bramREAD <= 0;
_q_uartInBuffer_wenable0 <= 0;
_q_uartInBuffer_addr0 <= 0;
_q_uartInBuffer_wenable1 <= 0;
_q_uartInBuffer_wdata1 <= 0;
_q_uartInBuffer_addr1 <= 0;
_q_uartInBufferNext <= 0;
_q_uartInBufferTop <= 0;
_q_uartInHold <= 1;
_q_uartOutBuffer_wenable0 <= 0;
_q_uartOutBuffer_addr0 <= 0;
_q_uartOutBuffer_wenable1 <= 0;
_q_uartOutBuffer_wdata1 <= 0;
_q_uartOutBuffer_addr1 <= 0;
_q_uartOutBufferNext <= 0;
_q_uartOutBufferTop <= 0;
_q_newuartOutBufferTop <= 0;
_q_uartOutHold <= 0;
  if (reset) begin
_q_index <= 0;
end else begin
_q_index <= 0;
end
  end else begin
_q_instruction <= _d_instruction;
_q_pc <= _d_pc;
_q_newPC <= _d_newPC;
_q_dstack_wenable <= _d_dstack_wenable;
_q_dstack_wdata <= _d_dstack_wdata;
_q_dstack_addr <= _d_dstack_addr;
_q_stackTop <= _d_stackTop;
_q_dsp <= _d_dsp;
_q_newDSP <= _d_newDSP;
_q_newStackTop <= _d_newStackTop;
_q_rstack_wenable <= _d_rstack_wenable;
_q_rstack_wdata <= _d_rstack_wdata;
_q_rstack_addr <= _d_rstack_addr;
_q_rsp <= _d_rsp;
_q_newRSP <= _d_newRSP;
_q_rstackWData <= _d_rstackWData;
_q_stackNext <= _d_stackNext;
_q_rStackTop <= _d_rStackTop;
_q_memoryInput <= _d_memoryInput;
_q_rom_addr <= _d_rom_addr;
_q_ram_wenable0 <= _d_ram_wenable0;
_q_ram_wdata0 <= _d_ram_wdata0;
_q_ram_addr0 <= _d_ram_addr0;
_q_ram_wenable1 <= _d_ram_wenable1;
_q_ram_addr1 <= _d_ram_addr1;
_q_CYCLE <= _d_CYCLE;
_q_INIT <= _d_INIT;
_q_copyaddress <= _d_copyaddress;
_q_bramREAD <= _d_bramREAD;
_q_uartInBuffer_wenable0 <= _d_uartInBuffer_wenable0;
_q_uartInBuffer_addr0 <= _d_uartInBuffer_addr0;
_q_uartInBuffer_wenable1 <= _d_uartInBuffer_wenable1;
_q_uartInBuffer_wdata1 <= _d_uartInBuffer_wdata1;
_q_uartInBuffer_addr1 <= _d_uartInBuffer_addr1;
_q_uartInBufferNext <= _d_uartInBufferNext;
_q_uartInBufferTop <= _d_uartInBufferTop;
_q_uartInHold <= _d_uartInHold;
_q_uartOutBuffer_wenable0 <= _d_uartOutBuffer_wenable0;
_q_uartOutBuffer_addr0 <= _d_uartOutBuffer_addr0;
_q_uartOutBuffer_wenable1 <= _d_uartOutBuffer_wenable1;
_q_uartOutBuffer_wdata1 <= _d_uartOutBuffer_wdata1;
_q_uartOutBuffer_addr1 <= _d_uartOutBuffer_addr1;
_q_uartOutBufferNext <= _d_uartOutBufferNext;
_q_uartOutBufferTop <= _d_uartOutBufferTop;
_q_newuartOutBufferTop <= _d_newuartOutBufferTop;
_q_uartOutHold <= _d_uartOutHold;
_q_index <= _d_index;
  end
_q_led <= _d_led;
_q_uart_tx_data <= _d_uart_tx_data;
_q_uart_tx_valid <= _d_uart_tx_valid;
_q_uart_rx_ready <= _d_uart_rx_ready;
_q_sdram_cle <= _d_sdram_cle;
_q_sdram_dqm <= _d_sdram_dqm;
_q_sdram_cs <= _d_sdram_cs;
_q_sdram_we <= _d_sdram_we;
_q_sdram_cas <= _d_sdram_cas;
_q_sdram_ras <= _d_sdram_ras;
_q_sdram_ba <= _d_sdram_ba;
_q_sdram_a <= _d_sdram_a;
_q_sdram_clk <= _d_sdram_clk;
_q_display_gpu_x <= _d_display_gpu_x;
_q_display_gpu_y <= _d_display_gpu_y;
_q_display_gpu_param0 <= _d_display_gpu_param0;
_q_display_gpu_param1 <= _d_display_gpu_param1;
_q_display_gpu_param2 <= _d_display_gpu_param2;
_q_display_gpu_param3 <= _d_display_gpu_param3;
_q_display_gpu_colour <= _d_display_gpu_colour;
_q_display_gpu_write <= _d_display_gpu_write;
_q_display_tpu_x <= _d_display_tpu_x;
_q_display_tpu_y <= _d_display_tpu_y;
_q_display_tpu_set <= _d_display_tpu_set;
_q_display_tpu_write <= _d_display_tpu_write;
_q_display_terminal_character <= _d_display_terminal_character;
_q_display_terminal_write <= _d_display_terminal_write;
_q_display_showterminal <= _d_display_showterminal;
_q_display_showcursor <= _d_display_showcursor;
end


reset_conditioner _vga_rstcond (
.rcclk(_w_clk_gen_outclk_1),
.in(reset),
.out(_w_vga_rstcond_out)
);

de10nano_clk_100_25 _clk_gen (
.refclk(clock),
.outclk_0(_w_clk_gen_outclk_0),
.outclk_1(_w_clk_gen_outclk_1),
.locked(_w_clk_gen_locked),
.rst(reset)
);
M_vga vga_driver (
.out_vga_hs(_w_vga_driver_vga_hs),
.out_vga_vs(_w_vga_driver_vga_vs),
.out_active(_w_vga_driver_active),
.out_vblank(_w_vga_driver_vblank),
.out_vga_x(_w_vga_driver_vga_x),
.out_vga_y(_w_vga_driver_vga_y),
.out_done(_w_vga_driver_done),
.in_run(_vga_driver_run),
.reset(_w_vga_rstcond_out),
.clock(_w_clk_gen_outclk_1)
);
M_multiplex_display display (
.in_pix_x(_w_vga_driver_vga_x),
.in_pix_y(_w_vga_driver_vga_y),
.in_pix_active(_w_vga_driver_active),
.in_pix_vblank(_w_vga_driver_vblank),
.in_gpu_x(_d_display_gpu_x),
.in_gpu_y(_d_display_gpu_y),
.in_gpu_param0(_d_display_gpu_param0),
.in_gpu_param1(_d_display_gpu_param1),
.in_gpu_param2(_d_display_gpu_param2),
.in_gpu_param3(_d_display_gpu_param3),
.in_gpu_colour(_d_display_gpu_colour),
.in_gpu_write(_d_display_gpu_write),
.in_tpu_x(_d_display_tpu_x),
.in_tpu_y(_d_display_tpu_y),
.in_tpu_set(_d_display_tpu_set),
.in_tpu_write(_d_display_tpu_write),
.in_terminal_character(_d_display_terminal_character),
.in_terminal_write(_d_display_terminal_write),
.in_showterminal(_d_display_showterminal),
.in_showcursor(_d_display_showcursor),
.in_timer1hz(in_timer1hz),
.out_pix_red(_w_display_pix_red),
.out_pix_green(_w_display_pix_green),
.out_pix_blue(_w_display_pix_blue),
.out_gpu_active(_w_display_gpu_active),
.out_done(_w_display_done),
.in_run(_display_run),
.reset(_w_vga_rstcond_out),
.clock(_w_clk_gen_outclk_1)
);

M_main_mem_dstack __mem__dstack(
.clock(clock),
.in_dstack_wenable(_d_dstack_wenable),
.in_dstack_wdata(_d_dstack_wdata),
.in_dstack_addr(_d_dstack_addr),
.out_dstack_rdata(_w_mem_dstack_rdata)
);
M_main_mem_rstack __mem__rstack(
.clock(clock),
.in_rstack_wenable(_d_rstack_wenable),
.in_rstack_wdata(_d_rstack_wdata),
.in_rstack_addr(_d_rstack_addr),
.out_rstack_rdata(_w_mem_rstack_rdata)
);
M_main_mem_rom __mem__rom(
.clock(clock),
.in_rom_addr(_d_rom_addr),
.out_rom_rdata(_w_mem_rom_rdata)
);
M_main_mem_ram __mem__ram(
.clock0(clock),
.clock1(clock),
.in_ram_wenable0(_d_ram_wenable0),
.in_ram_wdata0(_d_ram_wdata0),
.in_ram_addr0(_d_ram_addr0),
.in_ram_wenable1(_d_ram_wenable1),
.in_ram_wdata1(_c_ram_wdata1),
.in_ram_addr1(_d_ram_addr1),
.out_ram_rdata0(_w_mem_ram_rdata0),
.out_ram_rdata1(_w_mem_ram_rdata1)
);
M_main_mem_uartInBuffer __mem__uartInBuffer(
.clock0(clock),
.clock1(clock),
.in_uartInBuffer_wenable0(_d_uartInBuffer_wenable0),
.in_uartInBuffer_wdata0(_c_uartInBuffer_wdata0),
.in_uartInBuffer_addr0(_d_uartInBuffer_addr0),
.in_uartInBuffer_wenable1(_d_uartInBuffer_wenable1),
.in_uartInBuffer_wdata1(_d_uartInBuffer_wdata1),
.in_uartInBuffer_addr1(_d_uartInBuffer_addr1),
.out_uartInBuffer_rdata0(_w_mem_uartInBuffer_rdata0),
.out_uartInBuffer_rdata1(_w_mem_uartInBuffer_rdata1)
);
M_main_mem_uartOutBuffer __mem__uartOutBuffer(
.clock0(clock),
.clock1(clock),
.in_uartOutBuffer_wenable0(_d_uartOutBuffer_wenable0),
.in_uartOutBuffer_wdata0(_c_uartOutBuffer_wdata0),
.in_uartOutBuffer_addr0(_d_uartOutBuffer_addr0),
.in_uartOutBuffer_wenable1(_d_uartOutBuffer_wenable1),
.in_uartOutBuffer_wdata1(_d_uartOutBuffer_wdata1),
.in_uartOutBuffer_addr1(_d_uartOutBuffer_addr1),
.out_uartOutBuffer_rdata0(_w_mem_uartOutBuffer_rdata0),
.out_uartOutBuffer_rdata1(_w_mem_uartOutBuffer_rdata1)
);

assign _w_pcPlusOne = _d_pc+1;
assign _w_rdelta = {{7{_d_instruction[3+:1]}},_d_instruction[2+:1]};
assign _w_rstackWrite = (_w_is_call|(_w_is_alu&_d_instruction[6+:1]));
assign _w_dstackWrite = (_w_is_lit|(_w_is_alu&_d_instruction[7+:1]));
assign _w_ddelta = {{7{_d_instruction[1+:1]}},_d_instruction[0+:1]};
assign _w_is_call = (_d_instruction[13+:3]==3'b010);
assign _w_is_lit = _d_instruction[15+:1];
assign _w_is_alu = (_d_instruction[13+:3]==3'b011);
assign _w_immediate = (_d_instruction[0+:15]);

always @* begin
_d_instruction = _q_instruction;
_d_pc = _q_pc;
_d_newPC = _q_newPC;
_d_dstack_wenable = _q_dstack_wenable;
_d_dstack_wdata = _q_dstack_wdata;
_d_dstack_addr = _q_dstack_addr;
_d_stackTop = _q_stackTop;
_d_dsp = _q_dsp;
_d_newDSP = _q_newDSP;
_d_newStackTop = _q_newStackTop;
_d_rstack_wenable = _q_rstack_wenable;
_d_rstack_wdata = _q_rstack_wdata;
_d_rstack_addr = _q_rstack_addr;
_d_rsp = _q_rsp;
_d_newRSP = _q_newRSP;
_d_rstackWData = _q_rstackWData;
_d_stackNext = _q_stackNext;
_d_rStackTop = _q_rStackTop;
_d_memoryInput = _q_memoryInput;
_d_rom_addr = _q_rom_addr;
_d_ram_wenable0 = _q_ram_wenable0;
_d_ram_wdata0 = _q_ram_wdata0;
_d_ram_addr0 = _q_ram_addr0;
_d_ram_wenable1 = _q_ram_wenable1;
_d_ram_addr1 = _q_ram_addr1;
_d_CYCLE = _q_CYCLE;
_d_INIT = _q_INIT;
_d_copyaddress = _q_copyaddress;
_d_bramREAD = _q_bramREAD;
_d_uartInBuffer_wenable0 = _q_uartInBuffer_wenable0;
_d_uartInBuffer_addr0 = _q_uartInBuffer_addr0;
_d_uartInBuffer_wenable1 = _q_uartInBuffer_wenable1;
_d_uartInBuffer_wdata1 = _q_uartInBuffer_wdata1;
_d_uartInBuffer_addr1 = _q_uartInBuffer_addr1;
_d_uartInBufferNext = _q_uartInBufferNext;
_d_uartInBufferTop = _q_uartInBufferTop;
_d_uartInHold = _q_uartInHold;
_d_uartOutBuffer_wenable0 = _q_uartOutBuffer_wenable0;
_d_uartOutBuffer_addr0 = _q_uartOutBuffer_addr0;
_d_uartOutBuffer_wenable1 = _q_uartOutBuffer_wenable1;
_d_uartOutBuffer_wdata1 = _q_uartOutBuffer_wdata1;
_d_uartOutBuffer_addr1 = _q_uartOutBuffer_addr1;
_d_uartOutBufferNext = _q_uartOutBufferNext;
_d_uartOutBufferTop = _q_uartOutBufferTop;
_d_newuartOutBufferTop = _q_newuartOutBufferTop;
_d_uartOutHold = _q_uartOutHold;
_d_led = _q_led;
_d_uart_tx_data = _q_uart_tx_data;
_d_uart_tx_valid = _q_uart_tx_valid;
_d_uart_rx_ready = _q_uart_rx_ready;
_d_sdram_cle = _q_sdram_cle;
_d_sdram_dqm = _q_sdram_dqm;
_d_sdram_cs = _q_sdram_cs;
_d_sdram_we = _q_sdram_we;
_d_sdram_cas = _q_sdram_cas;
_d_sdram_ras = _q_sdram_ras;
_d_sdram_ba = _q_sdram_ba;
_d_sdram_a = _q_sdram_a;
_d_sdram_clk = _q_sdram_clk;
_d_display_gpu_x = _q_display_gpu_x;
_d_display_gpu_y = _q_display_gpu_y;
_d_display_gpu_param0 = _q_display_gpu_param0;
_d_display_gpu_param1 = _q_display_gpu_param1;
_d_display_gpu_param2 = _q_display_gpu_param2;
_d_display_gpu_param3 = _q_display_gpu_param3;
_d_display_gpu_colour = _q_display_gpu_colour;
_d_display_gpu_write = _q_display_gpu_write;
_d_display_tpu_x = _q_display_tpu_x;
_d_display_tpu_y = _q_display_tpu_y;
_d_display_tpu_set = _q_display_tpu_set;
_d_display_tpu_write = _q_display_tpu_write;
_d_display_terminal_character = _q_display_terminal_character;
_d_display_terminal_write = _q_display_terminal_write;
_d_display_showterminal = _q_display_showterminal;
_d_display_showcursor = _q_display_showcursor;
_d_index = _q_index;
_vga_driver_run = 1;
_display_run = 1;
// _always_pre
_d_dstack_wenable = 0;
_d_rstack_wenable = 0;
_d_uartInBuffer_wenable0 = 0;
_d_uartInBuffer_wenable1 = 1;
_d_uartInBuffer_addr0 = _q_uartInBufferNext;
_d_uartInBuffer_addr1 = _q_uartInBufferTop;
_d_uartOutBuffer_wenable0 = 0;
_d_uartOutBuffer_wenable1 = 1;
_d_uartOutBuffer_addr0 = _q_uartOutBufferNext;
_d_uartOutBuffer_addr1 = _q_uartOutBufferTop;
_d_sdram_cle = 1'bz;
_d_sdram_dqm = 1'bz;
_d_sdram_cs = 1'bz;
_d_sdram_we = 1'bz;
_d_sdram_cas = 1'bz;
_d_sdram_ras = 1'bz;
_d_sdram_ba = 2'bz;
_d_sdram_a = 13'bz;
_d_sdram_clk = 1'bz;
_d_index = 7;
case (_q_index)
0: begin
// _top
// var inits
_d_pc = 0;
_d_dstack_wenable = 0;
_d_dstack_wdata = 0;
_d_dstack_addr = 0;
_d_stackTop = 0;
_d_dsp = 0;
_d_rstack_wenable = 0;
_d_rstack_wdata = 0;
_d_rstack_addr = 0;
_d_rsp = 0;
_d_rom_addr = 0;
_d_ram_wenable0 = 0;
_d_ram_wdata0 = 0;
_d_ram_addr0 = 0;
_d_ram_wenable1 = 0;
_d_ram_addr1 = 0;
_d_CYCLE = 0;
_d_INIT = 0;
_d_copyaddress = 0;
_d_bramREAD = 0;
_d_uartInBuffer_wenable0 = 0;
_d_uartInBuffer_addr0 = 0;
_d_uartInBuffer_wenable1 = 0;
_d_uartInBuffer_wdata1 = 0;
_d_uartInBuffer_addr1 = 0;
_d_uartInBufferNext = 0;
_d_uartInBufferTop = 0;
_d_uartInHold = 1;
_d_uartOutBuffer_wenable0 = 0;
_d_uartOutBuffer_addr0 = 0;
_d_uartOutBuffer_wenable1 = 0;
_d_uartOutBuffer_wdata1 = 0;
_d_uartOutBuffer_addr1 = 0;
_d_uartOutBufferNext = 0;
_d_uartOutBufferTop = 0;
_d_newuartOutBufferTop = 0;
_d_uartOutHold = 0;
// --
_d_display_showterminal = 1;
_d_display_showcursor = 1;
_d_index = 1;
end
1: begin
// __while__block_1
if (_q_INIT==0) begin
// __block_2
// __block_4
  case (_q_CYCLE)
  0: begin
// __block_6_case
// __block_7
_d_ram_addr0 = _q_copyaddress;
_d_ram_wdata0 = 0;
_d_ram_wenable0 = 1;
// __block_8
  end
  1: begin
// __block_9_case
// __block_10
_d_copyaddress = _q_copyaddress+1;
_d_ram_wenable0 = 0;
// __block_11
  end
  4: begin
// __block_12_case
// __block_13
if (_q_copyaddress==32768) begin
// __block_14
// __block_16
_d_INIT = 1;
_d_copyaddress = 0;
// __block_17
end else begin
// __block_15
end
// __block_18
// __block_19
  end
  default: begin
// __block_20_case
// __block_21
// __block_22
  end
endcase
// __block_5
_d_CYCLE = (_q_CYCLE==4)?0:_q_CYCLE+1;
// __block_23
_d_index = 1;
end else begin
_d_index = 3;
end
end
3: begin
// __while__block_24
if (_q_INIT==1) begin
// __block_25
// __block_27
  case (_q_CYCLE)
  0: begin
// __block_29_case
// __block_30
_d_rom_addr = _q_copyaddress;
// __block_31
  end
  1: begin
// __block_32_case
// __block_33
_d_bramREAD = _w_mem_rom_rdata;
// __block_34
  end
  2: begin
// __block_35_case
// __block_36
_d_ram_addr0 = _q_copyaddress;
_d_ram_wdata0 = _q_bramREAD;
_d_ram_wenable0 = 1;
// __block_37
  end
  3: begin
// __block_38_case
// __block_39
_d_copyaddress = _q_copyaddress+1;
_d_ram_wenable0 = 0;
// __block_40
  end
  4: begin
// __block_41_case
// __block_42
if (_q_copyaddress==4096) begin
// __block_43
// __block_45
_d_INIT = 3;
_d_copyaddress = 0;
// __block_46
end else begin
// __block_44
end
// __block_47
// __block_48
  end
  default: begin
// __block_49_case
// __block_50
// __block_51
  end
endcase
// __block_28
_d_CYCLE = (_q_CYCLE==4)?0:_q_CYCLE+1;
// __block_52
_d_index = 3;
end else begin
_d_index = 5;
end
end
5: begin
// __while__block_53
if (_q_INIT==3) begin
// __block_54
// __block_56
  case (_q_uartInHold)
  0: begin
// __block_58_case
// __block_59
if (in_uart_rx_valid) begin
// __block_60
// __block_62
_d_uartInBuffer_wdata1 = in_uart_rx_data;
_d_uartInBufferTop = _q_uartInBufferTop+1;
_d_uartInHold = 1;
// __block_63
end else begin
// __block_61
end
// __block_64
_d_uart_rx_ready = 1;
// __block_65
  end
  1: begin
// __block_66_case
// __block_67
_d_uartInHold = (in_uart_rx_valid==0)?0:1;
// __block_68
  end
endcase
// __block_57
  case (_q_uartOutHold)
  0: begin
// __block_70_case
// __block_71
if (~(_q_uartOutBufferNext==_q_uartOutBufferTop)&~(in_uart_tx_busy)) begin
// __block_72
// __block_74
_d_uart_tx_data = _w_mem_uartOutBuffer_rdata0;
_d_uart_tx_valid = 1;
_d_uartOutHold = 1;
_d_uartOutBufferNext = _q_uartOutBufferNext+1;
// __block_75
end else begin
// __block_73
end
// __block_76
// __block_77
  end
  1: begin
// __block_78_case
// __block_79
if (~in_uart_tx_busy) begin
// __block_80
// __block_82
_d_uart_tx_valid = 0;
_d_uartOutHold = 0;
// __block_83
end else begin
// __block_81
end
// __block_84
// __block_85
  end
endcase
// __block_69
_d_uartOutBufferTop = _q_newuartOutBufferTop;
  case (_q_CYCLE)
  0: begin
// __block_87_case
// __block_88
_d_stackNext = _w_mem_dstack_rdata;
_d_rStackTop = _w_mem_rstack_rdata;
_d_ram_addr0 = _q_stackTop>>1;
_d_ram_wenable0 = 0;
_d_ram_addr1 = _q_pc;
_d_ram_wenable1 = 0;
// __block_89
  end
  1: begin
// __block_90_case
// __block_91
_d_memoryInput = _w_mem_ram_rdata0;
_d_instruction = _w_mem_ram_rdata1;
// __block_92
  end
  2: begin
// __block_93_case
// __block_94
if (_w_is_lit) begin
// __block_95
// __block_97
_d_newStackTop = _w_immediate;
_d_newPC = _w_pcPlusOne;
_d_newDSP = _q_dsp+1;
_d_newRSP = _q_rsp;
// __block_98
end else begin
// __block_96
// __block_99
  case (_q_instruction[13+:2])
  2'b00: begin
// __block_101_case
// __block_102
_d_newStackTop = _q_stackTop;
_d_newPC = _q_instruction[0+:13];
_d_newDSP = _q_dsp;
_d_newRSP = _q_rsp;
// __block_103
  end
  2'b01: begin
// __block_104_case
// __block_105
_d_newStackTop = _q_stackNext;
_d_newPC = (_q_stackTop==0)?_q_instruction[0+:13]:_w_pcPlusOne;
_d_newDSP = _q_dsp-1;
_d_newRSP = _q_rsp;
// __block_106
  end
  2'b10: begin
// __block_107_case
// __block_108
_d_newStackTop = _q_stackTop;
_d_newPC = _q_instruction[0+:13];
_d_newDSP = _q_dsp;
_d_newRSP = _q_rsp+1;
_d_rstackWData = _w_pcPlusOne<<1;
// __block_109
  end
  2'b11: begin
// __block_110_case
// __block_111
  case (_q_instruction[4+:1])
  1'b0: begin
// __block_113_case
// __block_114
  case (_q_instruction[8+:4])
  4'b0000: begin
// __block_116_case
// __block_117
_d_newStackTop = _q_stackTop;
// __block_118
  end
  4'b0001: begin
// __block_119_case
// __block_120
_d_newStackTop = _q_stackNext;
// __block_121
  end
  4'b0010: begin
// __block_122_case
// __block_123
_d_newStackTop = _q_stackTop+_q_stackNext;
// __block_124
  end
  4'b0011: begin
// __block_125_case
// __block_126
_d_newStackTop = _q_stackTop&_q_stackNext;
// __block_127
  end
  4'b0100: begin
// __block_128_case
// __block_129
_d_newStackTop = _q_stackTop|_q_stackNext;
// __block_130
  end
  4'b0101: begin
// __block_131_case
// __block_132
_d_newStackTop = _q_stackTop^_q_stackNext;
// __block_133
  end
  4'b0110: begin
// __block_134_case
// __block_135
_d_newStackTop = ~_q_stackTop;
// __block_136
  end
  4'b0111: begin
// __block_137_case
// __block_138
_d_newStackTop = {16{(_q_stackNext==_q_stackTop)}};
// __block_139
  end
  4'b1000: begin
// __block_140_case
// __block_141
_d_newStackTop = {16{($signed(_q_stackNext)<$signed(_q_stackTop))}};
// __block_142
  end
  4'b1001: begin
// __block_143_case
// __block_144
_d_newStackTop = _q_stackNext>>_q_stackTop[0+:4];
// __block_145
  end
  4'b1010: begin
// __block_146_case
// __block_147
_d_newStackTop = _q_stackTop-1;
// __block_148
  end
  4'b1011: begin
// __block_149_case
// __block_150
_d_newStackTop = _q_rStackTop;
// __block_151
  end
  4'b1100: begin
// __block_152_case
// __block_153
  case (_q_stackTop)
  16'hf000: begin
// __block_155_case
// __block_156
_d_newStackTop = {8'b0,_w_mem_uartInBuffer_rdata0};
_d_uartInBufferNext = _q_uartInBufferNext+1;
// __block_157
  end
  16'hf001: begin
// __block_158_case
// __block_159
_d_newStackTop = {14'b0,(_d_uartOutBufferTop+1==_d_uartOutBufferNext),~(_q_uartInBufferNext==_d_uartInBufferTop)};
// __block_160
  end
  16'hf002: begin
// __block_161_case
// __block_162
_d_newStackTop = _q_led;
// __block_163
  end
  16'hf003: begin
// __block_164_case
// __block_165
_d_newStackTop = {12'b0,in_buttons};
// __block_166
  end
  16'hf004: begin
// __block_167_case
// __block_168
_d_newStackTop = in_timer1hz;
// __block_169
  end
  16'hff07: begin
// __block_170_case
// __block_171
_d_newStackTop = _w_display_gpu_active;
// __block_172
  end
  default: begin
// __block_173_case
// __block_174
_d_newStackTop = _q_memoryInput;
// __block_175
  end
endcase
// __block_154
// __block_176
  end
  4'b1101: begin
// __block_177_case
// __block_178
_d_newStackTop = _q_stackNext<<_q_stackTop[0+:4];
// __block_179
  end
  4'b1110: begin
// __block_180_case
// __block_181
_d_newStackTop = {_q_rsp,_q_dsp};
// __block_182
  end
  4'b1111: begin
// __block_183_case
// __block_184
_d_newStackTop = {16{($unsigned(_q_stackNext)<$unsigned(_q_stackTop))}};
// __block_185
  end
endcase
// __block_115
// __block_186
  end
  1'b1: begin
// __block_187_case
// __block_188
  case (_q_instruction[8+:4])
  4'b0000: begin
// __block_190_case
// __block_191
_d_newStackTop = {16{(_q_stackTop==0)}};
// __block_192
  end
  4'b0001: begin
// __block_193_case
// __block_194
_d_newStackTop = ~{16{(_q_stackTop==0)}};
// __block_195
  end
  4'b0010: begin
// __block_196_case
// __block_197
_d_newStackTop = ~{16{(_q_stackNext==_q_stackTop)}};
// __block_198
  end
  4'b0011: begin
// __block_199_case
// __block_200
_d_newStackTop = _q_stackTop+1;
// __block_201
  end
  4'b0100: begin
// __block_202_case
// __block_203
_d_newStackTop = _q_stackTop<<1;
// __block_204
  end
  4'b0101: begin
// __block_205_case
// __block_206
_d_newStackTop = _q_stackTop>>1;
// __block_207
  end
  4'b0110: begin
// __block_208_case
// __block_209
_d_newStackTop = {16{($signed(_q_stackNext)>$signed(_q_stackTop))}};
// __block_210
  end
  4'b0111: begin
// __block_211_case
// __block_212
_d_newStackTop = {16{($unsigned(_q_stackNext)>$unsigned(_q_stackTop))}};
// __block_213
  end
  4'b1000: begin
// __block_214_case
// __block_215
_d_newStackTop = {16{($signed(_q_stackTop)<$signed(0))}};
// __block_216
  end
  4'b1001: begin
// __block_217_case
// __block_218
_d_newStackTop = {16{($signed(_q_stackTop)>$signed(0))}};
// __block_219
  end
  4'b1010: begin
// __block_220_case
// __block_221
_d_newStackTop = ($signed(_q_stackTop)<$signed(0))?-_q_stackTop:_q_stackTop;
// __block_222
  end
  4'b1011: begin
// __block_223_case
// __block_224
_d_newStackTop = ($signed(_q_stackNext)>$signed(_q_stackTop))?_q_stackNext:_q_stackTop;
// __block_225
  end
  4'b1100: begin
// __block_226_case
// __block_227
_d_newStackTop = ($signed(_q_stackNext)<$signed(_q_stackTop))?_q_stackNext:_q_stackTop;
// __block_228
  end
  4'b1101: begin
// __block_229_case
// __block_230
_d_newStackTop = -_q_stackTop;
// __block_231
  end
  4'b1110: begin
// __block_232_case
// __block_233
_d_newStackTop = _q_stackNext-_q_stackTop;
// __block_234
  end
  4'b1111: begin
// __block_235_case
// __block_236
_d_newStackTop = {16{($signed(_q_stackNext)>=$signed(_q_stackTop))}};
// __block_237
  end
endcase
// __block_189
// __block_238
  end
endcase
// __block_112
_d_newDSP = _q_dsp+_w_ddelta;
_d_newRSP = _q_rsp+_w_rdelta;
_d_rstackWData = _q_stackTop;
_d_newPC = (_q_instruction[12+:1])?_q_rStackTop>>1:_w_pcPlusOne;
if (_q_instruction[5+:1]) begin
// __block_239
// __block_241
  case (_q_stackTop)
  default: begin
// __block_243_case
// __block_244
_d_ram_addr0 = _q_stackTop>>1;
_d_ram_wdata0 = _q_stackNext;
_d_ram_wenable0 = 1;
// __block_245
  end
  16'hf000: begin
// __block_246_case
// __block_247
_d_uartOutBuffer_wdata1 = _q_stackNext[0+:8];
_d_newuartOutBufferTop = _d_uartOutBufferTop+1;
// __block_248
  end
  16'hf002: begin
// __block_249_case
// __block_250
_d_led = _q_stackNext;
// __block_251
  end
  16'hff00: begin
// __block_252_case
// __block_253
_d_display_gpu_x = _q_stackNext;
// __block_254
  end
  16'hff01: begin
// __block_255_case
// __block_256
_d_display_gpu_y = _q_stackNext;
// __block_257
  end
  16'hff02: begin
// __block_258_case
// __block_259
_d_display_gpu_colour = _q_stackNext;
// __block_260
  end
  16'hff03: begin
// __block_261_case
// __block_262
_d_display_gpu_param0 = _q_stackNext;
// __block_263
  end
  16'hff04: begin
// __block_264_case
// __block_265
_d_display_gpu_param1 = _q_stackNext;
// __block_266
  end
  16'hff05: begin
// __block_267_case
// __block_268
_d_display_gpu_param2 = _q_stackNext;
// __block_269
  end
  16'hff06: begin
// __block_270_case
// __block_271
_d_display_gpu_param3 = _q_stackNext;
// __block_272
  end
  16'hff07: begin
// __block_273_case
// __block_274
_d_display_gpu_write = _q_stackNext;
// __block_275
  end
  16'hff10: begin
// __block_276_case
// __block_277
_d_display_tpu_x = _q_stackNext;
// __block_278
  end
  16'hff11: begin
// __block_279_case
// __block_280
_d_display_tpu_y = _q_stackNext;
// __block_281
  end
  16'hff12: begin
// __block_282_case
// __block_283
_d_display_tpu_set = _q_stackNext;
_d_display_tpu_write = 1;
// __block_284
  end
  16'hff13: begin
// __block_285_case
// __block_286
_d_display_tpu_set = _q_stackNext;
_d_display_tpu_write = 2;
// __block_287
  end
  16'hff14: begin
// __block_288_case
// __block_289
_d_display_tpu_set = _q_stackNext;
_d_display_tpu_write = 3;
// __block_290
  end
  16'hff20: begin
// __block_291_case
// __block_292
_d_display_terminal_character = _q_stackNext;
_d_display_terminal_write = 1;
// __block_293
  end
  16'hff21: begin
// __block_294_case
// __block_295
_d_display_showterminal = _q_stackNext;
// __block_296
  end
endcase
// __block_242
// __block_297
end else begin
// __block_240
end
// __block_298
// __block_299
  end
endcase
// __block_100
// __block_300
end
// __block_301
// __block_302
  end
  3: begin
// __block_303_case
// __block_304
if (_w_dstackWrite) begin
// __block_305
// __block_307
_d_dstack_wenable = 1;
_d_dstack_addr = _q_newDSP;
_d_dstack_wdata = _q_stackTop;
// __block_308
end else begin
// __block_306
end
// __block_309
if (_w_rstackWrite) begin
// __block_310
// __block_312
_d_rstack_wenable = 1;
_d_rstack_addr = _q_newRSP;
_d_rstack_wdata = _q_rstackWData;
// __block_313
end else begin
// __block_311
end
// __block_314
// __block_315
  end
  4: begin
// __block_316_case
// __block_317
_d_dsp = _q_newDSP;
_d_pc = _q_newPC;
_d_stackTop = _q_newStackTop;
_d_rsp = _q_newRSP;
_d_dstack_addr = _q_newDSP;
_d_rstack_addr = _q_newRSP;
_d_ram_wenable0 = 0;
_d_display_gpu_write = 0;
_d_display_tpu_write = 0;
_d_display_terminal_write = 0;
// __block_318
  end
  default: begin
// __block_319_case
// __block_320
// __block_321
  end
endcase
// __block_86
_d_CYCLE = (_q_CYCLE==4)?0:_q_CYCLE+1;
// __block_322
_d_index = 5;
end else begin
_d_index = 6;
end
end
6: begin
// __block_55
_d_index = 7;
end
7: begin // end of main
end
default: begin 
_d_index = 7;
 end
endcase
end
endmodule

